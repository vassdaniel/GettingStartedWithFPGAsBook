// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 27 2024 21:36:36

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "State_Machine_Top" view "INTERFACE"

module State_Machine_Top (
    o_Segment2_D,
    o_LED_3,
    i_Switch_4,
    i_Clk,
    o_Segment2_G,
    o_Segment2_C,
    o_LED_2,
    i_Switch_1,
    o_Segment2_F,
    o_Segment2_B,
    o_LED_1,
    i_Switch_2,
    o_Segment2_E,
    o_Segment2_A,
    o_LED_4,
    i_Switch_3);

    output o_Segment2_D;
    output o_LED_3;
    input i_Switch_4;
    input i_Clk;
    output o_Segment2_G;
    output o_Segment2_C;
    output o_LED_2;
    input i_Switch_1;
    output o_Segment2_F;
    output o_Segment2_B;
    output o_LED_1;
    input i_Switch_2;
    output o_Segment2_E;
    output o_Segment2_A;
    output o_LED_4;
    input i_Switch_3;

    wire N__8507;
    wire N__8506;
    wire N__8505;
    wire N__8496;
    wire N__8495;
    wire N__8494;
    wire N__8487;
    wire N__8486;
    wire N__8485;
    wire N__8478;
    wire N__8477;
    wire N__8476;
    wire N__8469;
    wire N__8468;
    wire N__8467;
    wire N__8460;
    wire N__8459;
    wire N__8458;
    wire N__8451;
    wire N__8450;
    wire N__8449;
    wire N__8442;
    wire N__8441;
    wire N__8440;
    wire N__8433;
    wire N__8432;
    wire N__8431;
    wire N__8424;
    wire N__8423;
    wire N__8422;
    wire N__8415;
    wire N__8414;
    wire N__8413;
    wire N__8406;
    wire N__8405;
    wire N__8404;
    wire N__8397;
    wire N__8396;
    wire N__8395;
    wire N__8388;
    wire N__8387;
    wire N__8386;
    wire N__8379;
    wire N__8378;
    wire N__8377;
    wire N__8370;
    wire N__8369;
    wire N__8368;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8332;
    wire N__8331;
    wire N__8328;
    wire N__8325;
    wire N__8322;
    wire N__8319;
    wire N__8314;
    wire N__8313;
    wire N__8308;
    wire N__8305;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8287;
    wire N__8286;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8267;
    wire N__8266;
    wire N__8265;
    wire N__8264;
    wire N__8263;
    wire N__8262;
    wire N__8261;
    wire N__8260;
    wire N__8259;
    wire N__8258;
    wire N__8257;
    wire N__8256;
    wire N__8255;
    wire N__8254;
    wire N__8253;
    wire N__8252;
    wire N__8251;
    wire N__8250;
    wire N__8249;
    wire N__8248;
    wire N__8247;
    wire N__8246;
    wire N__8245;
    wire N__8244;
    wire N__8243;
    wire N__8242;
    wire N__8241;
    wire N__8240;
    wire N__8239;
    wire N__8238;
    wire N__8237;
    wire N__8236;
    wire N__8235;
    wire N__8234;
    wire N__8233;
    wire N__8232;
    wire N__8231;
    wire N__8230;
    wire N__8229;
    wire N__8228;
    wire N__8227;
    wire N__8226;
    wire N__8225;
    wire N__8224;
    wire N__8223;
    wire N__8222;
    wire N__8221;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8119;
    wire N__8118;
    wire N__8117;
    wire N__8110;
    wire N__8107;
    wire N__8102;
    wire N__8101;
    wire N__8098;
    wire N__8095;
    wire N__8092;
    wire N__8089;
    wire N__8084;
    wire N__8083;
    wire N__8082;
    wire N__8075;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8062;
    wire N__8057;
    wire N__8056;
    wire N__8053;
    wire N__8052;
    wire N__8051;
    wire N__8048;
    wire N__8047;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8037;
    wire N__8034;
    wire N__8031;
    wire N__8028;
    wire N__8027;
    wire N__8024;
    wire N__8017;
    wire N__8016;
    wire N__8011;
    wire N__8008;
    wire N__8003;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7985;
    wire N__7982;
    wire N__7981;
    wire N__7980;
    wire N__7979;
    wire N__7976;
    wire N__7971;
    wire N__7968;
    wire N__7961;
    wire N__7960;
    wire N__7957;
    wire N__7954;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7936;
    wire N__7935;
    wire N__7934;
    wire N__7931;
    wire N__7926;
    wire N__7923;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7885;
    wire N__7882;
    wire N__7877;
    wire N__7874;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7853;
    wire N__7852;
    wire N__7849;
    wire N__7846;
    wire N__7845;
    wire N__7844;
    wire N__7843;
    wire N__7832;
    wire N__7831;
    wire N__7830;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7816;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7802;
    wire N__7801;
    wire N__7798;
    wire N__7793;
    wire N__7792;
    wire N__7787;
    wire N__7782;
    wire N__7779;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7765;
    wire N__7764;
    wire N__7763;
    wire N__7762;
    wire N__7761;
    wire N__7750;
    wire N__7747;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7737;
    wire N__7736;
    wire N__7731;
    wire N__7730;
    wire N__7727;
    wire N__7724;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7712;
    wire N__7709;
    wire N__7700;
    wire N__7699;
    wire N__7698;
    wire N__7697;
    wire N__7696;
    wire N__7693;
    wire N__7690;
    wire N__7687;
    wire N__7686;
    wire N__7681;
    wire N__7680;
    wire N__7679;
    wire N__7676;
    wire N__7671;
    wire N__7668;
    wire N__7665;
    wire N__7660;
    wire N__7659;
    wire N__7658;
    wire N__7657;
    wire N__7656;
    wire N__7655;
    wire N__7654;
    wire N__7653;
    wire N__7652;
    wire N__7645;
    wire N__7642;
    wire N__7639;
    wire N__7632;
    wire N__7625;
    wire N__7620;
    wire N__7617;
    wire N__7604;
    wire N__7603;
    wire N__7602;
    wire N__7601;
    wire N__7600;
    wire N__7599;
    wire N__7596;
    wire N__7595;
    wire N__7594;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7576;
    wire N__7573;
    wire N__7568;
    wire N__7567;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7559;
    wire N__7558;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7544;
    wire N__7541;
    wire N__7540;
    wire N__7535;
    wire N__7528;
    wire N__7525;
    wire N__7522;
    wire N__7519;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7503;
    wire N__7484;
    wire N__7483;
    wire N__7480;
    wire N__7479;
    wire N__7476;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7468;
    wire N__7467;
    wire N__7464;
    wire N__7461;
    wire N__7460;
    wire N__7455;
    wire N__7452;
    wire N__7449;
    wire N__7446;
    wire N__7443;
    wire N__7440;
    wire N__7437;
    wire N__7434;
    wire N__7431;
    wire N__7418;
    wire N__7417;
    wire N__7416;
    wire N__7415;
    wire N__7414;
    wire N__7413;
    wire N__7410;
    wire N__7407;
    wire N__7406;
    wire N__7405;
    wire N__7404;
    wire N__7403;
    wire N__7402;
    wire N__7399;
    wire N__7398;
    wire N__7397;
    wire N__7394;
    wire N__7393;
    wire N__7388;
    wire N__7387;
    wire N__7386;
    wire N__7381;
    wire N__7376;
    wire N__7369;
    wire N__7364;
    wire N__7361;
    wire N__7356;
    wire N__7353;
    wire N__7348;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7322;
    wire N__7319;
    wire N__7316;
    wire N__7315;
    wire N__7314;
    wire N__7313;
    wire N__7310;
    wire N__7303;
    wire N__7300;
    wire N__7299;
    wire N__7296;
    wire N__7293;
    wire N__7290;
    wire N__7283;
    wire N__7282;
    wire N__7281;
    wire N__7278;
    wire N__7277;
    wire N__7270;
    wire N__7267;
    wire N__7262;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7252;
    wire N__7251;
    wire N__7250;
    wire N__7249;
    wire N__7238;
    wire N__7237;
    wire N__7236;
    wire N__7235;
    wire N__7234;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7219;
    wire N__7214;
    wire N__7211;
    wire N__7210;
    wire N__7207;
    wire N__7204;
    wire N__7199;
    wire N__7196;
    wire N__7187;
    wire N__7186;
    wire N__7183;
    wire N__7180;
    wire N__7175;
    wire N__7174;
    wire N__7171;
    wire N__7168;
    wire N__7165;
    wire N__7160;
    wire N__7157;
    wire N__7156;
    wire N__7153;
    wire N__7150;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7136;
    wire N__7133;
    wire N__7130;
    wire N__7127;
    wire N__7124;
    wire N__7121;
    wire N__7118;
    wire N__7115;
    wire N__7114;
    wire N__7113;
    wire N__7112;
    wire N__7109;
    wire N__7106;
    wire N__7105;
    wire N__7102;
    wire N__7099;
    wire N__7098;
    wire N__7095;
    wire N__7094;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7071;
    wire N__7066;
    wire N__7061;
    wire N__7052;
    wire N__7049;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7039;
    wire N__7036;
    wire N__7033;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7021;
    wire N__7018;
    wire N__7015;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7003;
    wire N__7000;
    wire N__6997;
    wire N__6992;
    wire N__6991;
    wire N__6988;
    wire N__6985;
    wire N__6980;
    wire N__6977;
    wire N__6974;
    wire N__6971;
    wire N__6970;
    wire N__6969;
    wire N__6968;
    wire N__6967;
    wire N__6964;
    wire N__6961;
    wire N__6958;
    wire N__6957;
    wire N__6956;
    wire N__6945;
    wire N__6942;
    wire N__6939;
    wire N__6938;
    wire N__6935;
    wire N__6932;
    wire N__6929;
    wire N__6928;
    wire N__6925;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6902;
    wire N__6899;
    wire N__6892;
    wire N__6889;
    wire N__6884;
    wire N__6881;
    wire N__6880;
    wire N__6877;
    wire N__6874;
    wire N__6871;
    wire N__6866;
    wire N__6865;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6852;
    wire N__6845;
    wire N__6842;
    wire N__6841;
    wire N__6838;
    wire N__6835;
    wire N__6830;
    wire N__6827;
    wire N__6826;
    wire N__6823;
    wire N__6820;
    wire N__6815;
    wire N__6812;
    wire N__6811;
    wire N__6808;
    wire N__6805;
    wire N__6800;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6790;
    wire N__6787;
    wire N__6784;
    wire N__6781;
    wire N__6776;
    wire N__6775;
    wire N__6774;
    wire N__6773;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6755;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6727;
    wire N__6724;
    wire N__6721;
    wire N__6716;
    wire N__6713;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6701;
    wire N__6698;
    wire N__6697;
    wire N__6694;
    wire N__6691;
    wire N__6686;
    wire N__6683;
    wire N__6682;
    wire N__6681;
    wire N__6678;
    wire N__6673;
    wire N__6668;
    wire N__6665;
    wire N__6664;
    wire N__6661;
    wire N__6658;
    wire N__6653;
    wire N__6650;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6638;
    wire N__6635;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6625;
    wire N__6620;
    wire N__6617;
    wire N__6616;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6602;
    wire N__6599;
    wire N__6598;
    wire N__6597;
    wire N__6594;
    wire N__6589;
    wire N__6584;
    wire N__6581;
    wire N__6580;
    wire N__6579;
    wire N__6576;
    wire N__6571;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6557;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6545;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6530;
    wire N__6529;
    wire N__6524;
    wire N__6521;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6509;
    wire N__6508;
    wire N__6505;
    wire N__6502;
    wire N__6497;
    wire N__6496;
    wire N__6493;
    wire N__6490;
    wire N__6487;
    wire N__6482;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6470;
    wire N__6469;
    wire N__6464;
    wire N__6461;
    wire N__6458;
    wire N__6457;
    wire N__6454;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6437;
    wire N__6436;
    wire N__6435;
    wire N__6432;
    wire N__6431;
    wire N__6426;
    wire N__6423;
    wire N__6420;
    wire N__6413;
    wire N__6412;
    wire N__6411;
    wire N__6410;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6394;
    wire N__6393;
    wire N__6392;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6374;
    wire N__6373;
    wire N__6370;
    wire N__6369;
    wire N__6366;
    wire N__6363;
    wire N__6360;
    wire N__6353;
    wire N__6352;
    wire N__6349;
    wire N__6346;
    wire N__6341;
    wire N__6338;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6305;
    wire N__6302;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6290;
    wire N__6287;
    wire N__6286;
    wire N__6283;
    wire N__6280;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6248;
    wire N__6247;
    wire N__6244;
    wire N__6241;
    wire N__6236;
    wire N__6235;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6221;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6209;
    wire N__6208;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6188;
    wire N__6187;
    wire N__6186;
    wire N__6183;
    wire N__6178;
    wire N__6173;
    wire N__6170;
    wire N__6169;
    wire N__6164;
    wire N__6161;
    wire N__6160;
    wire N__6157;
    wire N__6154;
    wire N__6149;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6137;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6125;
    wire N__6122;
    wire N__6119;
    wire N__6116;
    wire N__6113;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6086;
    wire N__6083;
    wire N__6080;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6067;
    wire N__6066;
    wire N__6063;
    wire N__6060;
    wire N__6057;
    wire N__6052;
    wire N__6049;
    wire N__6044;
    wire N__6043;
    wire N__6042;
    wire N__6037;
    wire N__6034;
    wire N__6029;
    wire N__6026;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6014;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__5999;
    wire N__5998;
    wire N__5995;
    wire N__5992;
    wire N__5987;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5947;
    wire N__5944;
    wire N__5941;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5900;
    wire N__5899;
    wire N__5896;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5886;
    wire N__5879;
    wire N__5878;
    wire N__5877;
    wire N__5874;
    wire N__5873;
    wire N__5868;
    wire N__5865;
    wire N__5862;
    wire N__5855;
    wire N__5854;
    wire N__5853;
    wire N__5852;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5813;
    wire N__5812;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5802;
    wire N__5799;
    wire N__5796;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5782;
    wire N__5781;
    wire N__5778;
    wire N__5775;
    wire N__5772;
    wire N__5767;
    wire N__5762;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5754;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5729;
    wire N__5728;
    wire N__5725;
    wire N__5722;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5710;
    wire N__5707;
    wire N__5704;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5683;
    wire N__5682;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5665;
    wire N__5662;
    wire N__5661;
    wire N__5658;
    wire N__5657;
    wire N__5652;
    wire N__5649;
    wire N__5648;
    wire N__5647;
    wire N__5644;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5634;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5620;
    wire N__5617;
    wire N__5612;
    wire N__5603;
    wire N__5602;
    wire N__5601;
    wire N__5594;
    wire N__5593;
    wire N__5592;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5554;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5542;
    wire N__5537;
    wire N__5534;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5522;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5486;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5474;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5459;
    wire N__5456;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5434;
    wire N__5431;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5416;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5390;
    wire N__5387;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5364;
    wire N__5363;
    wire N__5358;
    wire N__5353;
    wire N__5348;
    wire N__5345;
    wire N__5344;
    wire N__5341;
    wire N__5340;
    wire N__5339;
    wire N__5338;
    wire N__5337;
    wire N__5336;
    wire N__5335;
    wire N__5334;
    wire N__5333;
    wire N__5332;
    wire N__5331;
    wire N__5330;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5314;
    wire N__5305;
    wire N__5300;
    wire N__5297;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5252;
    wire N__5249;
    wire N__5248;
    wire N__5247;
    wire N__5246;
    wire N__5245;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5231;
    wire N__5228;
    wire N__5219;
    wire N__5216;
    wire N__5215;
    wire N__5214;
    wire N__5213;
    wire N__5212;
    wire N__5211;
    wire N__5208;
    wire N__5201;
    wire N__5196;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5167;
    wire N__5166;
    wire N__5163;
    wire N__5158;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5098;
    wire N__5097;
    wire N__5090;
    wire N__5087;
    wire N__5086;
    wire N__5083;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5068;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5054;
    wire N__5051;
    wire N__5048;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5033;
    wire N__5030;
    wire N__5029;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5014;
    wire N__5009;
    wire N__5006;
    wire N__5005;
    wire N__5002;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4987;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4966;
    wire N__4965;
    wire N__4964;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4945;
    wire N__4942;
    wire N__4939;
    wire N__4936;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4924;
    wire N__4921;
    wire N__4918;
    wire N__4915;
    wire N__4910;
    wire N__4909;
    wire N__4906;
    wire N__4903;
    wire N__4898;
    wire N__4895;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4880;
    wire N__4877;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4865;
    wire N__4862;
    wire N__4861;
    wire N__4858;
    wire N__4855;
    wire N__4850;
    wire N__4847;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4835;
    wire N__4832;
    wire N__4831;
    wire N__4830;
    wire N__4827;
    wire N__4822;
    wire N__4817;
    wire N__4814;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4802;
    wire N__4799;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4750;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4732;
    wire N__4731;
    wire N__4730;
    wire N__4725;
    wire N__4722;
    wire N__4719;
    wire N__4712;
    wire N__4711;
    wire N__4708;
    wire N__4707;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4691;
    wire N__4688;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4669;
    wire N__4668;
    wire N__4665;
    wire N__4664;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4646;
    wire N__4643;
    wire N__4642;
    wire N__4639;
    wire N__4636;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4603;
    wire N__4600;
    wire N__4599;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4587;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4570;
    wire N__4569;
    wire N__4568;
    wire N__4563;
    wire N__4558;
    wire N__4553;
    wire N__4550;
    wire N__4549;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4504;
    wire N__4503;
    wire N__4500;
    wire N__4495;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4483;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4459;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4445;
    wire N__4442;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4430;
    wire N__4427;
    wire N__4426;
    wire N__4423;
    wire N__4420;
    wire N__4417;
    wire N__4412;
    wire N__4409;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4397;
    wire N__4394;
    wire N__4393;
    wire N__4390;
    wire N__4387;
    wire N__4382;
    wire N__4379;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4367;
    wire N__4364;
    wire N__4363;
    wire N__4360;
    wire N__4357;
    wire N__4352;
    wire N__4349;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4334;
    wire N__4331;
    wire N__4330;
    wire N__4329;
    wire N__4328;
    wire N__4327;
    wire N__4326;
    wire N__4325;
    wire N__4324;
    wire N__4323;
    wire N__4322;
    wire N__4321;
    wire N__4320;
    wire N__4319;
    wire N__4310;
    wire N__4307;
    wire N__4302;
    wire N__4299;
    wire N__4294;
    wire N__4287;
    wire N__4282;
    wire N__4271;
    wire N__4268;
    wire N__4267;
    wire N__4264;
    wire N__4261;
    wire N__4258;
    wire N__4253;
    wire N__4252;
    wire N__4251;
    wire N__4250;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4223;
    wire N__4220;
    wire N__4219;
    wire N__4216;
    wire N__4213;
    wire N__4208;
    wire N__4205;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4190;
    wire N__4187;
    wire N__4186;
    wire N__4183;
    wire N__4180;
    wire N__4175;
    wire N__4172;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4160;
    wire N__4157;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4145;
    wire N__4142;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4127;
    wire N__4124;
    wire N__4123;
    wire N__4120;
    wire N__4117;
    wire N__4112;
    wire N__4109;
    wire N__4108;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4084;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4074;
    wire N__4067;
    wire N__4066;
    wire N__4065;
    wire N__4062;
    wire N__4061;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4043;
    wire N__4042;
    wire N__4039;
    wire N__4036;
    wire N__4031;
    wire N__4028;
    wire N__4027;
    wire N__4024;
    wire N__4021;
    wire N__4016;
    wire N__4013;
    wire N__4010;
    wire N__4009;
    wire N__4006;
    wire N__4003;
    wire N__4000;
    wire N__3995;
    wire N__3992;
    wire N__3991;
    wire N__3988;
    wire N__3985;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3953;
    wire N__3950;
    wire N__3949;
    wire N__3946;
    wire N__3943;
    wire N__3938;
    wire N__3935;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3923;
    wire N__3922;
    wire N__3919;
    wire N__3916;
    wire N__3911;
    wire N__3910;
    wire N__3907;
    wire N__3904;
    wire N__3899;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3887;
    wire N__3886;
    wire N__3883;
    wire N__3880;
    wire N__3875;
    wire N__3874;
    wire N__3871;
    wire N__3868;
    wire N__3863;
    wire N__3862;
    wire N__3859;
    wire N__3856;
    wire N__3851;
    wire N__3848;
    wire N__3847;
    wire N__3844;
    wire N__3841;
    wire N__3838;
    wire N__3833;
    wire N__3832;
    wire N__3829;
    wire N__3826;
    wire N__3821;
    wire N__3818;
    wire N__3815;
    wire N__3812;
    wire N__3809;
    wire N__3806;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3794;
    wire N__3791;
    wire N__3788;
    wire N__3787;
    wire N__3784;
    wire N__3781;
    wire N__3776;
    wire N__3775;
    wire N__3772;
    wire N__3769;
    wire N__3764;
    wire N__3763;
    wire N__3760;
    wire N__3757;
    wire N__3754;
    wire N__3749;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3680;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3668;
    wire N__3665;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3629;
    wire N__3626;
    wire GNDG0;
    wire VCCG0;
    wire bfn_4_7_0_;
    wire \Debounce_SW1.un2_r_count_cry_1 ;
    wire \Debounce_SW1.un2_r_count_cry_2 ;
    wire \Debounce_SW1.un2_r_count_cry_3 ;
    wire \Debounce_SW1.un2_r_count_cry_4 ;
    wire \Debounce_SW1.un2_r_count_cry_5 ;
    wire \Debounce_SW1.un2_r_count_cry_6 ;
    wire \Debounce_SW1.un2_r_count_cry_7 ;
    wire \Debounce_SW1.un2_r_count_cry_8 ;
    wire bfn_4_8_0_;
    wire \Debounce_SW1.un2_r_count_cry_9 ;
    wire \Debounce_SW1.un2_r_count_cry_10 ;
    wire \Debounce_SW1.un2_r_count_cry_11 ;
    wire \Debounce_SW1.un2_r_count_cry_12 ;
    wire \Debounce_SW1.un2_r_count_cry_13 ;
    wire \Debounce_SW1.un2_r_count_cry_14 ;
    wire \Debounce_SW1.un2_r_count_cry_15 ;
    wire \Debounce_SW1.un2_r_count_cry_16 ;
    wire bfn_4_9_0_;
    wire \Game_Inst.N_83_i ;
    wire r_Hex_Encoding_i_1;
    wire r_Hex_Encoding_i_4;
    wire r_Hex_Encoding_i_5;
    wire r_Hex_Encoding_i_6;
    wire r_Hex_Encoding_i_0;
    wire r_Hex_Encoding_i_3;
    wire \Game_Inst.Count_Inst.un4_i_enable_12_cascade_ ;
    wire \Debounce_SW1.r_CountZ0Z_6 ;
    wire \Debounce_SW1.r_CountZ0Z_5 ;
    wire \Debounce_SW1.r_CountZ0Z_4 ;
    wire \Debounce_SW1.r_CountZ0Z_16 ;
    wire \Debounce_SW1.r_CountZ0Z_15 ;
    wire \Debounce_SW1.r_CountZ0Z_17 ;
    wire \Debounce_SW1.r_CountZ0Z_14 ;
    wire \Game_Inst.Count_Inst.un4_i_enable_16_cascade_ ;
    wire \Game_Inst.Count_Inst.un4_i_enable_8 ;
    wire \Game_Inst.Count_Inst.un4_i_enable_17 ;
    wire \Game_Inst.Count_Inst.un4_i_enable_14 ;
    wire \Game_Inst.Count_Inst.un4_i_enable_19_cascade_ ;
    wire \Game_Inst.Count_Inst.un4_i_enable_13 ;
    wire \Debounce_SW1.r_CountZ0Z_10 ;
    wire \Debounce_SW1.r_CountZ0Z_9 ;
    wire \Debounce_SW1.r_CountZ0Z_11 ;
    wire \Debounce_SW1.r_CountZ0Z_8 ;
    wire \Game_Inst.r_SM_Main_ns_i_0_a2_0_0_0_cascade_ ;
    wire \Game_Inst.N_346 ;
    wire \Game_Inst.N_346_cascade_ ;
    wire \Game_Inst.o_Toggle_4_i_43 ;
    wire \Game_Inst.LFSR_Inst.r_LFSRZ0Z_16 ;
    wire \Game_Inst.LFSR_Inst.r_LFSRZ0Z_17 ;
    wire \Game_Inst.LFSR_Inst.r_LFSRZ0Z_18 ;
    wire \Game_Inst.LFSR_Inst.r_LFSRZ0Z_19 ;
    wire \Game_Inst.w_LFSR_Data_0 ;
    wire \Game_Inst.LFSR_Inst.r_LFSRZ0Z_20 ;
    wire \Game_Inst.LFSR_Inst.r_LFSRZ0Z_21 ;
    wire r_Hex_Encoding_i_2;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_1 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_0 ;
    wire bfn_6_6_0_;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_2 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_1 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_3 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_2 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_4 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_3 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_5 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_4 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_6 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_5 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_7 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_6 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_8 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_7 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_8 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_9 ;
    wire bfn_6_7_0_;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_10 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_9 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_11 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_10 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_12 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_11 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_13 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_12 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_14 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_13 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_15 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_14 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_16 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_15 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_16 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_17 ;
    wire bfn_6_8_0_;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_18 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_17 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_19 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_18 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_20 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_19 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_21 ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_20 ;
    wire \Game_Inst.Count_Inst.un4_i_enable ;
    wire \Game_Inst.Count_Inst.un2_r_counter_cry_21 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_22 ;
    wire \Game_Inst.N_83_i_g ;
    wire \Game_Inst.N_128_cascade_ ;
    wire \Game_Inst.N_130 ;
    wire \Game_Inst.N_130_cascade_ ;
    wire \Game_Inst.r_Index_0_sqmuxa_2_i_2_0 ;
    wire \Game_Inst.r_Index_0_sqmuxa_2_i_1_0_cascade_ ;
    wire \Game_Inst.N_209_cascade_ ;
    wire \Game_Inst.N_91_2 ;
    wire \Game_Inst.N_210_cascade_ ;
    wire \Game_Inst.SUM_i_i_0_1 ;
    wire \Game_Inst.r_Pattern_0Z0Z_0 ;
    wire \Game_Inst.r_Pattern_1Z0Z_0 ;
    wire \Game_Inst.r_Pattern_0_RNIDQ911Z0Z_0_cascade_ ;
    wire \Game_Inst.un6_r_button_dv_7_i_m2_ns_1_0_cascade_ ;
    wire \Game_Inst.N_145 ;
    wire \Game_Inst.SUM_i_i_0_tz_0 ;
    wire \Game_Inst.N_91 ;
    wire \Game_Inst.r_SM_Main_ns_i_i_o2_0_1_1_cascade_ ;
    wire \Game_Inst.r_Pattern_7Z0Z_0 ;
    wire \Game_Inst.r_Pattern_6Z0Z_0 ;
    wire \Game_Inst.r_Pattern_6_RNIPUEEZ0Z_0 ;
    wire \Game_Inst.N_132 ;
    wire \Game_Inst.N_132_cascade_ ;
    wire \Game_Inst.w_LFSR_Data_14 ;
    wire \Game_Inst.N_262 ;
    wire \Game_Inst.r_SM_Main_ns_i_i_a2_1_0_1 ;
    wire \Game_Inst.r_SM_Main_ns_i_i_1_1_cascade_ ;
    wire \Game_Inst.r_SM_Main_ns_i_i_3_1_cascade_ ;
    wire \Game_Inst.N_137 ;
    wire \Game_Inst.N_128 ;
    wire \Debounce_SW4.N_181_cascade_ ;
    wire \Debounce_SW4.N_42 ;
    wire \Debounce_SW4.un9_r_count_10_cascade_ ;
    wire \Debounce_SW4.N_288 ;
    wire \Debounce_SW4.N_158 ;
    wire \Debounce_SW4.N_158_cascade_ ;
    wire \Debounce_SW4.N_149 ;
    wire \Debounce_SW4.un9_r_count_10 ;
    wire \Debounce_SW4.un9_r_count_0_a2_2_cascade_ ;
    wire \Debounce_SW4.r_CountZ0Z_0 ;
    wire \Debounce_SW4.r_CountZ0Z_1 ;
    wire bfn_7_5_0_;
    wire \Debounce_SW4.r_CountZ0Z_2 ;
    wire \Debounce_SW4.un2_r_count_cry_1 ;
    wire \Debounce_SW4.r_CountZ0Z_3 ;
    wire \Debounce_SW4.un2_r_count_cry_2 ;
    wire \Debounce_SW4.r_CountZ0Z_4 ;
    wire \Debounce_SW4.un2_r_count_cry_3 ;
    wire \Debounce_SW4.r_CountZ0Z_5 ;
    wire \Debounce_SW4.un2_r_count_cry_4 ;
    wire \Debounce_SW4.r_CountZ0Z_6 ;
    wire \Debounce_SW4.un2_r_count_cry_5 ;
    wire \Debounce_SW4.r_CountZ0Z_7 ;
    wire \Debounce_SW4.un2_r_count_cry_6 ;
    wire \Debounce_SW4.r_CountZ0Z_8 ;
    wire \Debounce_SW4.un2_r_count_cry_7 ;
    wire \Debounce_SW4.un2_r_count_cry_8 ;
    wire \Debounce_SW4.r_CountZ0Z_9 ;
    wire bfn_7_6_0_;
    wire \Debounce_SW4.r_CountZ0Z_10 ;
    wire \Debounce_SW4.un2_r_count_cry_9 ;
    wire \Debounce_SW4.r_CountZ0Z_11 ;
    wire \Debounce_SW4.un2_r_count_cry_10 ;
    wire \Debounce_SW4.r_CountZ0Z_12 ;
    wire \Debounce_SW4.un2_r_count_cry_11 ;
    wire \Debounce_SW4.r_CountZ0Z_13 ;
    wire \Debounce_SW4.un2_r_count_cry_12 ;
    wire \Debounce_SW4.un2_r_count_cry_13 ;
    wire \Debounce_SW4.un2_r_count_cry_14 ;
    wire \Debounce_SW4.un2_r_count_cry_15 ;
    wire \Debounce_SW4.un2_r_count_cry_16 ;
    wire bfn_7_7_0_;
    wire \Debounce_SW4.N_42_g ;
    wire \Debounce_SW1.r_CountZ0Z_2 ;
    wire \Debounce_SW1.r_CountZ0Z_3 ;
    wire \Debounce_SW1.un9_r_count_10_cascade_ ;
    wire \Debounce_SW1.N_285_cascade_ ;
    wire \Debounce_SW1.N_184_cascade_ ;
    wire \Debounce_SW1.N_36 ;
    wire \Game_Inst.r_Button_IDZ0Z_0 ;
    wire \Game_Inst.N_255_cascade_ ;
    wire \Game_Inst.N_167 ;
    wire \Game_Inst.N_255 ;
    wire \Game_Inst.r_Button_IDZ0Z_1 ;
    wire \Game_Inst.r_IndexZ0Z_1 ;
    wire \Game_Inst.r_Pattern_0_RNIFS911Z0Z_1_cascade_ ;
    wire \Game_Inst.r_IndexZ0Z_2 ;
    wire \Game_Inst.un6_r_button_dv_7_i_m2_ns_1_1_cascade_ ;
    wire \Game_Inst.r_Pattern_3_RNIH6MLZ0Z_0 ;
    wire \Game_Inst.r_Pattern_3_RNIJ8MLZ0Z_1 ;
    wire \Game_Inst.N_303 ;
    wire \Game_Inst.r_SM_Main_ns_i_0_2_0 ;
    wire \Game_Inst.r_Pattern_6_RNIR0FEZ0Z_1 ;
    wire \Game_Inst.r_Pattern_4_RNINK2AZ0Z_1 ;
    wire \Game_Inst.N_266 ;
    wire \Game_Inst.r_Button_DVZ0 ;
    wire \Game_Inst.r_SM_Main_d_6_cascade_ ;
    wire \Game_Inst.r_IndexZ1Z_0 ;
    wire \Game_Inst.r_Pattern_4_RNILI2AZ0Z_0 ;
    wire \Game_Inst.N_259 ;
    wire \Game_Inst.r_SM_Main_ns_i_0_1_2_cascade_ ;
    wire \Game_Inst.N_260_1 ;
    wire bfn_7_13_0_;
    wire \Debounce_SW2.un2_r_count_cry_1 ;
    wire \Debounce_SW2.un2_r_count_cry_2 ;
    wire \Debounce_SW2.un2_r_count_cry_3 ;
    wire \Debounce_SW2.un2_r_count_cry_4 ;
    wire \Debounce_SW2.un2_r_count_cry_5 ;
    wire \Debounce_SW2.un2_r_count_cry_6 ;
    wire \Debounce_SW2.un2_r_count_cry_7 ;
    wire \Debounce_SW2.un2_r_count_cry_8 ;
    wire bfn_7_14_0_;
    wire \Debounce_SW2.un2_r_count_cry_9 ;
    wire \Debounce_SW2.un2_r_count_cry_10 ;
    wire \Debounce_SW2.un2_r_count_cry_11 ;
    wire \Debounce_SW2.un2_r_count_cry_12 ;
    wire \Debounce_SW2.un2_r_count_cry_13 ;
    wire \Debounce_SW2.un2_r_count_cry_14 ;
    wire \Debounce_SW2.un2_r_count_cry_15 ;
    wire \Debounce_SW2.un2_r_count_cry_16 ;
    wire bfn_7_15_0_;
    wire i_Switch_4_c;
    wire \Debounce_SW4.r_State_e_0_RNO_2 ;
    wire \Debounce_SW3.N_159 ;
    wire \Debounce_SW3.N_159_cascade_ ;
    wire \Debounce_SW3.N_287 ;
    wire \Debounce_SW3.un9_r_count_0_a2_2 ;
    wire \Debounce_SW3.N_148 ;
    wire \Debounce_SW3.r_count15_i_a2_0_cascade_ ;
    wire \Debounce_SW3.un9_r_count_10 ;
    wire \Debounce_SW4.r_CountZ0Z_15 ;
    wire \Debounce_SW4.r_CountZ0Z_16 ;
    wire \Debounce_SW4.r_CountZ0Z_14 ;
    wire \Debounce_SW4.r_CountZ0Z_17 ;
    wire \Debounce_SW4.r_count15_i_a2_0 ;
    wire \Debounce_SW1.r_CountZ0Z_1 ;
    wire \Debounce_SW1.r_CountZ0Z_0 ;
    wire \Debounce_SW1.N_36_g ;
    wire \Debounce_SW1.N_146 ;
    wire \Debounce_SW1.r_CountZ0Z_12 ;
    wire \Debounce_SW1.r_CountZ0Z_13 ;
    wire \Debounce_SW1.r_CountZ0Z_7 ;
    wire \Debounce_SW1.un9_r_count_10 ;
    wire \Debounce_SW1.r_count15_i_a2_0 ;
    wire \Debounce_SW1.un9_r_count_0_a2_2_cascade_ ;
    wire \Debounce_SW1.N_161 ;
    wire \Game_Inst.r_SwitchZ0Z_4 ;
    wire \Game_Inst.r_SwitchZ0Z_2 ;
    wire \Game_Inst.r_Switch_1_RNIA12HZ0 ;
    wire \Game_Inst.r_SwitchZ0Z_1 ;
    wire \Game_Inst.w_Toggle ;
    wire \Game_Inst.r_ToggleZ0 ;
    wire \Game_Inst.N_208_cascade_ ;
    wire \Game_Inst.N_264 ;
    wire \Game_Inst.r_Pattern_5Z0Z_0 ;
    wire \Game_Inst.r_Pattern_3Z0Z_1 ;
    wire \Game_Inst.r_Pattern_2Z0Z_1 ;
    wire \Game_Inst.w_LFSR_Data_1 ;
    wire \Game_Inst.r_Pattern_0Z0Z_1 ;
    wire \Game_Inst.r_Pattern_1Z0Z_1 ;
    wire \Game_Inst.r_Pattern_6Z0Z_1 ;
    wire \Game_Inst.r_Pattern_2Z0Z_0 ;
    wire \Game_Inst.r_Pattern_3Z0Z_0 ;
    wire \Game_Inst.r_Pattern_4Z0Z_1 ;
    wire \Game_Inst.r_Pattern_4Z0Z_0 ;
    wire \Game_Inst.w_LFSR_Data_15 ;
    wire \Game_Inst.r_Pattern_7Z0Z_1 ;
    wire \Game_Inst.r_Pattern_5Z0Z_1 ;
    wire \Game_Inst.r_SM_Main_d_6 ;
    wire N_143;
    wire \Game_Inst.w_LFSR_Data_7 ;
    wire \Game_Inst.w_LFSR_Data_2 ;
    wire \Game_Inst.w_LFSR_Data_6 ;
    wire \Game_Inst.w_LFSR_Data_5 ;
    wire \Game_Inst.w_LFSR_Data_3 ;
    wire \Game_Inst.w_LFSR_Data_4 ;
    wire \Debounce_SW2.N_183_cascade_ ;
    wire \Debounce_SW2.N_38 ;
    wire \Debounce_SW2.r_CountZ0Z_10 ;
    wire \Debounce_SW2.r_CountZ0Z_9 ;
    wire \Debounce_SW2.r_CountZ0Z_11 ;
    wire \Debounce_SW2.r_CountZ0Z_8 ;
    wire \Debounce_SW2.r_CountZ0Z_13 ;
    wire \Debounce_SW2.r_CountZ0Z_12 ;
    wire \Debounce_SW2.un9_r_count_0_a2_2_cascade_ ;
    wire \Debounce_SW2.N_160 ;
    wire \Debounce_SW2.r_CountZ0Z_6 ;
    wire \Debounce_SW2.r_CountZ0Z_5 ;
    wire \Debounce_SW2.r_CountZ0Z_4 ;
    wire \Debounce_SW2.N_147 ;
    wire \Debounce_SW2.r_CountZ0Z_7 ;
    wire \Debounce_SW2.N_147_cascade_ ;
    wire \Debounce_SW2.N_286 ;
    wire \Debounce_SW2.r_CountZ0Z_2 ;
    wire \Debounce_SW2.r_CountZ0Z_3 ;
    wire \Debounce_SW2.un9_r_count_10 ;
    wire \Debounce_SW2.r_CountZ0Z_16 ;
    wire \Debounce_SW2.r_CountZ0Z_15 ;
    wire \Debounce_SW2.r_CountZ0Z_17 ;
    wire \Debounce_SW2.r_CountZ0Z_14 ;
    wire \Debounce_SW2.r_count15_i_a2_0 ;
    wire \Debounce_SW2.r_CountZ0Z_1 ;
    wire \Debounce_SW2.r_CountZ0Z_0 ;
    wire \Debounce_SW2.N_38_g ;
    wire \Debounce_SW3.r_CountZ0Z_0 ;
    wire \Debounce_SW3.r_CountZ0Z_1 ;
    wire bfn_9_5_0_;
    wire \Debounce_SW3.r_CountZ0Z_2 ;
    wire \Debounce_SW3.un2_r_count_cry_1 ;
    wire \Debounce_SW3.r_CountZ0Z_3 ;
    wire \Debounce_SW3.un2_r_count_cry_2 ;
    wire \Debounce_SW3.r_CountZ0Z_4 ;
    wire \Debounce_SW3.un2_r_count_cry_3 ;
    wire \Debounce_SW3.r_CountZ0Z_5 ;
    wire \Debounce_SW3.un2_r_count_cry_4 ;
    wire \Debounce_SW3.r_CountZ0Z_6 ;
    wire \Debounce_SW3.un2_r_count_cry_5 ;
    wire \Debounce_SW3.r_CountZ0Z_7 ;
    wire \Debounce_SW3.un2_r_count_cry_6 ;
    wire \Debounce_SW3.r_CountZ0Z_8 ;
    wire \Debounce_SW3.un2_r_count_cry_7 ;
    wire \Debounce_SW3.un2_r_count_cry_8 ;
    wire \Debounce_SW3.r_CountZ0Z_9 ;
    wire bfn_9_6_0_;
    wire \Debounce_SW3.r_CountZ0Z_10 ;
    wire \Debounce_SW3.un2_r_count_cry_9 ;
    wire \Debounce_SW3.r_CountZ0Z_11 ;
    wire \Debounce_SW3.un2_r_count_cry_10 ;
    wire \Debounce_SW3.r_CountZ0Z_12 ;
    wire \Debounce_SW3.un2_r_count_cry_11 ;
    wire \Debounce_SW3.r_CountZ0Z_13 ;
    wire \Debounce_SW3.un2_r_count_cry_12 ;
    wire \Debounce_SW3.r_CountZ0Z_14 ;
    wire \Debounce_SW3.un2_r_count_cry_13 ;
    wire \Debounce_SW3.r_CountZ0Z_15 ;
    wire \Debounce_SW3.un2_r_count_cry_14 ;
    wire \Debounce_SW3.r_CountZ0Z_16 ;
    wire \Debounce_SW3.un2_r_count_cry_15 ;
    wire \Debounce_SW3.un2_r_count_cry_16 ;
    wire bfn_9_7_0_;
    wire \Debounce_SW3.r_CountZ0Z_17 ;
    wire \Debounce_SW3.N_40_g ;
    wire i_Switch_1_c;
    wire \Debounce_SW1.r_State_e_0_RNOZ0 ;
    wire \Game_Inst.w_LFSR_Data_11 ;
    wire \Game_Inst.w_LFSR_Data_12 ;
    wire \Game_Inst.w_LFSR_Data_13 ;
    wire \Game_Inst.w_LFSR_Data_10 ;
    wire bfn_9_11_0_;
    wire \Game_Inst.un1_r_Score_cry_0 ;
    wire \Game_Inst.un1_r_Score_cry_1 ;
    wire \Game_Inst.un1_r_Score_cry_2 ;
    wire w_Score_3;
    wire \Game_Inst.N_291_cascade_ ;
    wire \Game_Inst.N_68_i ;
    wire \Game_Inst.un1_r_Score_cry_0_THRU_CO ;
    wire w_Score_1;
    wire \Game_Inst.r_Score_RNO_0Z0Z_0 ;
    wire w_Score_0;
    wire \Game_Inst.r_SM_MainZ0Z_0 ;
    wire \Game_Inst.r_SM_MainZ0Z_2 ;
    wire \Game_Inst.N_291 ;
    wire \Game_Inst.r_SM_MainZ0Z_1 ;
    wire \Game_Inst.N_241 ;
    wire \Game_Inst.r_Score_0_sqmuxa ;
    wire \Game_Inst.un1_r_SM_Main_0 ;
    wire \Game_Inst.N_241_cascade_ ;
    wire \Game_Inst.r_Score_RNO_0Z0Z_2 ;
    wire w_Score_2;
    wire \Game_Inst.w_LFSR_Data_8 ;
    wire \Game_Inst.w_LFSR_Data_9 ;
    wire i_Switch_2_c;
    wire \Debounce_SW2.r_State_e_0_RNOZ0Z_0 ;
    wire \Debounce_SW3.r_State_e_0_RNO_1 ;
    wire w_Switch_1;
    wire N_70;
    wire N_44;
    wire w_Switch_4;
    wire N_89;
    wire \Game_Inst.N_140 ;
    wire \Game_Inst.r_SwitchZ0Z_3 ;
    wire i_Clk_c_g;
    wire \Game_Inst.N_17 ;
    wire \Game_Inst.N_338 ;
    wire w_Switch_2;
    wire \Game_Inst.N_16 ;
    wire N_87;
    wire w_Switch_3;
    wire \Debounce_SW3.r_count15_i_a2_0 ;
    wire i_Switch_3_c;
    wire \Debounce_SW3.N_182 ;
    wire \Debounce_SW3.N_40 ;
    wire _gnd_net_;

    PRE_IO_GBUF i_Clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__8505),
            .GLOBALBUFFEROUTPUT(i_Clk_c_g));
    IO_PAD i_Clk_ibuf_gb_io_iopad (
            .OE(N__8507),
            .DIN(N__8506),
            .DOUT(N__8505),
            .PACKAGEPIN(i_Clk));
    defparam i_Clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam i_Clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Clk_ibuf_gb_io_preio (
            .PADOEN(N__8507),
            .PADOUT(N__8506),
            .PADIN(N__8505),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_F_obuf_iopad (
            .OE(N__8496),
            .DIN(N__8495),
            .DOUT(N__8494),
            .PACKAGEPIN(o_Segment2_F));
    defparam o_Segment2_F_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_F_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_F_obuf_preio (
            .PADOEN(N__8496),
            .PADOUT(N__8495),
            .PADIN(N__8494),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3659),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_1_obuf_iopad (
            .OE(N__8487),
            .DIN(N__8486),
            .DOUT(N__8485),
            .PACKAGEPIN(o_LED_1));
    defparam o_LED_1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_1_obuf_preio (
            .PADOEN(N__8487),
            .PADOUT(N__8486),
            .PADIN(N__8485),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7052),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_4_ibuf_iopad (
            .OE(N__8478),
            .DIN(N__8477),
            .DOUT(N__8476),
            .PACKAGEPIN(i_Switch_4));
    defparam i_Switch_4_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_4_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_4_ibuf_preio (
            .PADOEN(N__8478),
            .PADOUT(N__8477),
            .PADIN(N__8476),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_4_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_1_ibuf_iopad (
            .OE(N__8469),
            .DIN(N__8468),
            .DOUT(N__8467),
            .PACKAGEPIN(i_Switch_1));
    defparam i_Switch_1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_1_ibuf_preio (
            .PADOEN(N__8469),
            .PADOUT(N__8468),
            .PADIN(N__8467),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_3_ibuf_iopad (
            .OE(N__8460),
            .DIN(N__8459),
            .DOUT(N__8458),
            .PACKAGEPIN(i_Switch_3));
    defparam i_Switch_3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_3_ibuf_preio (
            .PADOEN(N__8460),
            .PADOUT(N__8459),
            .PADIN(N__8458),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_2_obuf_iopad (
            .OE(N__8451),
            .DIN(N__8450),
            .DOUT(N__8449),
            .PACKAGEPIN(o_LED_2));
    defparam o_LED_2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_2_obuf_preio (
            .PADOEN(N__8451),
            .PADOUT(N__8450),
            .PADIN(N__8449),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7949),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_E_obuf_iopad (
            .OE(N__8442),
            .DIN(N__8441),
            .DOUT(N__8440),
            .PACKAGEPIN(o_Segment2_E));
    defparam o_Segment2_E_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_E_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_E_obuf_preio (
            .PADOEN(N__8442),
            .PADOUT(N__8441),
            .PADIN(N__8440),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4094),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_C_obuf_iopad (
            .OE(N__8433),
            .DIN(N__8432),
            .DOUT(N__8431),
            .PACKAGEPIN(o_Segment2_C));
    defparam o_Segment2_C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_C_obuf_preio (
            .PADOEN(N__8433),
            .PADOUT(N__8432),
            .PADIN(N__8431),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3737),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_4_obuf_iopad (
            .OE(N__8424),
            .DIN(N__8423),
            .DOUT(N__8422),
            .PACKAGEPIN(o_LED_4));
    defparam o_LED_4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_4_obuf_preio (
            .PADOEN(N__8424),
            .PADOUT(N__8423),
            .PADIN(N__8422),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8300),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_B_obuf_iopad (
            .OE(N__8415),
            .DIN(N__8414),
            .DOUT(N__8413),
            .PACKAGEPIN(o_Segment2_B));
    defparam o_Segment2_B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_B_obuf_preio (
            .PADOEN(N__8415),
            .PADOUT(N__8414),
            .PADIN(N__8413),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3731),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_3_obuf_iopad (
            .OE(N__8406),
            .DIN(N__8405),
            .DOUT(N__8404),
            .PACKAGEPIN(o_LED_3));
    defparam o_LED_3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_3_obuf_preio (
            .PADOEN(N__8406),
            .PADOUT(N__8405),
            .PADIN(N__8404),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8351),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_A_obuf_iopad (
            .OE(N__8397),
            .DIN(N__8396),
            .DOUT(N__8395),
            .PACKAGEPIN(o_Segment2_A));
    defparam o_Segment2_A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_A_obuf_preio (
            .PADOEN(N__8397),
            .PADOUT(N__8396),
            .PADIN(N__8395),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3719),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_G_obuf_iopad (
            .OE(N__8388),
            .DIN(N__8387),
            .DOUT(N__8386),
            .PACKAGEPIN(o_Segment2_G));
    defparam o_Segment2_G_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_G_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_G_obuf_preio (
            .PADOEN(N__8388),
            .PADOUT(N__8387),
            .PADIN(N__8386),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3707),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_D_obuf_iopad (
            .OE(N__8379),
            .DIN(N__8378),
            .DOUT(N__8377),
            .PACKAGEPIN(o_Segment2_D));
    defparam o_Segment2_D_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_D_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_D_obuf_preio (
            .PADOEN(N__8379),
            .PADOUT(N__8378),
            .PADIN(N__8377),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3701),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_2_ibuf_iopad (
            .OE(N__8370),
            .DIN(N__8369),
            .DOUT(N__8368),
            .PACKAGEPIN(i_Switch_2));
    defparam i_Switch_2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_2_ibuf_preio (
            .PADOEN(N__8370),
            .PADOUT(N__8369),
            .PADIN(N__8368),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__1888 (
            .O(N__8351),
            .I(N__8348));
    LocalMux I__1887 (
            .O(N__8348),
            .I(N__8345));
    Span4Mux_s1_h I__1886 (
            .O(N__8345),
            .I(N__8342));
    Odrv4 I__1885 (
            .O(N__8342),
            .I(N_44));
    CascadeMux I__1884 (
            .O(N__8339),
            .I(N__8336));
    InMux I__1883 (
            .O(N__8336),
            .I(N__8333));
    LocalMux I__1882 (
            .O(N__8333),
            .I(N__8328));
    InMux I__1881 (
            .O(N__8332),
            .I(N__8325));
    InMux I__1880 (
            .O(N__8331),
            .I(N__8322));
    Span4Mux_v I__1879 (
            .O(N__8328),
            .I(N__8319));
    LocalMux I__1878 (
            .O(N__8325),
            .I(N__8314));
    LocalMux I__1877 (
            .O(N__8322),
            .I(N__8314));
    Span4Mux_h I__1876 (
            .O(N__8319),
            .I(N__8308));
    Span4Mux_v I__1875 (
            .O(N__8314),
            .I(N__8308));
    InMux I__1874 (
            .O(N__8313),
            .I(N__8305));
    Odrv4 I__1873 (
            .O(N__8308),
            .I(w_Switch_4));
    LocalMux I__1872 (
            .O(N__8305),
            .I(w_Switch_4));
    IoInMux I__1871 (
            .O(N__8300),
            .I(N__8297));
    LocalMux I__1870 (
            .O(N__8297),
            .I(N__8294));
    Odrv4 I__1869 (
            .O(N__8294),
            .I(N_89));
    CascadeMux I__1868 (
            .O(N__8291),
            .I(N__8288));
    InMux I__1867 (
            .O(N__8288),
            .I(N__8279));
    InMux I__1866 (
            .O(N__8287),
            .I(N__8279));
    InMux I__1865 (
            .O(N__8286),
            .I(N__8279));
    LocalMux I__1864 (
            .O(N__8279),
            .I(N__8276));
    Odrv12 I__1863 (
            .O(N__8276),
            .I(\Game_Inst.N_140 ));
    InMux I__1862 (
            .O(N__8273),
            .I(N__8270));
    LocalMux I__1861 (
            .O(N__8270),
            .I(\Game_Inst.r_SwitchZ0Z_3 ));
    ClkMux I__1860 (
            .O(N__8267),
            .I(N__8126));
    ClkMux I__1859 (
            .O(N__8266),
            .I(N__8126));
    ClkMux I__1858 (
            .O(N__8265),
            .I(N__8126));
    ClkMux I__1857 (
            .O(N__8264),
            .I(N__8126));
    ClkMux I__1856 (
            .O(N__8263),
            .I(N__8126));
    ClkMux I__1855 (
            .O(N__8262),
            .I(N__8126));
    ClkMux I__1854 (
            .O(N__8261),
            .I(N__8126));
    ClkMux I__1853 (
            .O(N__8260),
            .I(N__8126));
    ClkMux I__1852 (
            .O(N__8259),
            .I(N__8126));
    ClkMux I__1851 (
            .O(N__8258),
            .I(N__8126));
    ClkMux I__1850 (
            .O(N__8257),
            .I(N__8126));
    ClkMux I__1849 (
            .O(N__8256),
            .I(N__8126));
    ClkMux I__1848 (
            .O(N__8255),
            .I(N__8126));
    ClkMux I__1847 (
            .O(N__8254),
            .I(N__8126));
    ClkMux I__1846 (
            .O(N__8253),
            .I(N__8126));
    ClkMux I__1845 (
            .O(N__8252),
            .I(N__8126));
    ClkMux I__1844 (
            .O(N__8251),
            .I(N__8126));
    ClkMux I__1843 (
            .O(N__8250),
            .I(N__8126));
    ClkMux I__1842 (
            .O(N__8249),
            .I(N__8126));
    ClkMux I__1841 (
            .O(N__8248),
            .I(N__8126));
    ClkMux I__1840 (
            .O(N__8247),
            .I(N__8126));
    ClkMux I__1839 (
            .O(N__8246),
            .I(N__8126));
    ClkMux I__1838 (
            .O(N__8245),
            .I(N__8126));
    ClkMux I__1837 (
            .O(N__8244),
            .I(N__8126));
    ClkMux I__1836 (
            .O(N__8243),
            .I(N__8126));
    ClkMux I__1835 (
            .O(N__8242),
            .I(N__8126));
    ClkMux I__1834 (
            .O(N__8241),
            .I(N__8126));
    ClkMux I__1833 (
            .O(N__8240),
            .I(N__8126));
    ClkMux I__1832 (
            .O(N__8239),
            .I(N__8126));
    ClkMux I__1831 (
            .O(N__8238),
            .I(N__8126));
    ClkMux I__1830 (
            .O(N__8237),
            .I(N__8126));
    ClkMux I__1829 (
            .O(N__8236),
            .I(N__8126));
    ClkMux I__1828 (
            .O(N__8235),
            .I(N__8126));
    ClkMux I__1827 (
            .O(N__8234),
            .I(N__8126));
    ClkMux I__1826 (
            .O(N__8233),
            .I(N__8126));
    ClkMux I__1825 (
            .O(N__8232),
            .I(N__8126));
    ClkMux I__1824 (
            .O(N__8231),
            .I(N__8126));
    ClkMux I__1823 (
            .O(N__8230),
            .I(N__8126));
    ClkMux I__1822 (
            .O(N__8229),
            .I(N__8126));
    ClkMux I__1821 (
            .O(N__8228),
            .I(N__8126));
    ClkMux I__1820 (
            .O(N__8227),
            .I(N__8126));
    ClkMux I__1819 (
            .O(N__8226),
            .I(N__8126));
    ClkMux I__1818 (
            .O(N__8225),
            .I(N__8126));
    ClkMux I__1817 (
            .O(N__8224),
            .I(N__8126));
    ClkMux I__1816 (
            .O(N__8223),
            .I(N__8126));
    ClkMux I__1815 (
            .O(N__8222),
            .I(N__8126));
    ClkMux I__1814 (
            .O(N__8221),
            .I(N__8126));
    GlobalMux I__1813 (
            .O(N__8126),
            .I(N__8123));
    gio2CtrlBuf I__1812 (
            .O(N__8123),
            .I(i_Clk_c_g));
    InMux I__1811 (
            .O(N__8120),
            .I(N__8110));
    InMux I__1810 (
            .O(N__8119),
            .I(N__8110));
    InMux I__1809 (
            .O(N__8118),
            .I(N__8110));
    InMux I__1808 (
            .O(N__8117),
            .I(N__8107));
    LocalMux I__1807 (
            .O(N__8110),
            .I(N__8102));
    LocalMux I__1806 (
            .O(N__8107),
            .I(N__8102));
    Span4Mux_v I__1805 (
            .O(N__8102),
            .I(N__8098));
    CascadeMux I__1804 (
            .O(N__8101),
            .I(N__8095));
    Sp12to4 I__1803 (
            .O(N__8098),
            .I(N__8092));
    InMux I__1802 (
            .O(N__8095),
            .I(N__8089));
    Odrv12 I__1801 (
            .O(N__8092),
            .I(\Game_Inst.N_17 ));
    LocalMux I__1800 (
            .O(N__8089),
            .I(\Game_Inst.N_17 ));
    InMux I__1799 (
            .O(N__8084),
            .I(N__8075));
    InMux I__1798 (
            .O(N__8083),
            .I(N__8075));
    InMux I__1797 (
            .O(N__8082),
            .I(N__8075));
    LocalMux I__1796 (
            .O(N__8075),
            .I(N__8071));
    InMux I__1795 (
            .O(N__8074),
            .I(N__8068));
    Span4Mux_v I__1794 (
            .O(N__8071),
            .I(N__8065));
    LocalMux I__1793 (
            .O(N__8068),
            .I(N__8062));
    Odrv4 I__1792 (
            .O(N__8065),
            .I(\Game_Inst.N_338 ));
    Odrv12 I__1791 (
            .O(N__8062),
            .I(\Game_Inst.N_338 ));
    CascadeMux I__1790 (
            .O(N__8057),
            .I(N__8053));
    CascadeMux I__1789 (
            .O(N__8056),
            .I(N__8048));
    InMux I__1788 (
            .O(N__8053),
            .I(N__8043));
    InMux I__1787 (
            .O(N__8052),
            .I(N__8040));
    InMux I__1786 (
            .O(N__8051),
            .I(N__8037));
    InMux I__1785 (
            .O(N__8048),
            .I(N__8034));
    InMux I__1784 (
            .O(N__8047),
            .I(N__8031));
    InMux I__1783 (
            .O(N__8046),
            .I(N__8028));
    LocalMux I__1782 (
            .O(N__8043),
            .I(N__8024));
    LocalMux I__1781 (
            .O(N__8040),
            .I(N__8017));
    LocalMux I__1780 (
            .O(N__8037),
            .I(N__8017));
    LocalMux I__1779 (
            .O(N__8034),
            .I(N__8017));
    LocalMux I__1778 (
            .O(N__8031),
            .I(N__8011));
    LocalMux I__1777 (
            .O(N__8028),
            .I(N__8011));
    InMux I__1776 (
            .O(N__8027),
            .I(N__8008));
    Span4Mux_s3_h I__1775 (
            .O(N__8024),
            .I(N__8003));
    Span4Mux_h I__1774 (
            .O(N__8017),
            .I(N__8003));
    InMux I__1773 (
            .O(N__8016),
            .I(N__8000));
    Span4Mux_h I__1772 (
            .O(N__8011),
            .I(N__7997));
    LocalMux I__1771 (
            .O(N__8008),
            .I(N__7994));
    Odrv4 I__1770 (
            .O(N__8003),
            .I(w_Switch_2));
    LocalMux I__1769 (
            .O(N__8000),
            .I(w_Switch_2));
    Odrv4 I__1768 (
            .O(N__7997),
            .I(w_Switch_2));
    Odrv4 I__1767 (
            .O(N__7994),
            .I(w_Switch_2));
    CascadeMux I__1766 (
            .O(N__7985),
            .I(N__7982));
    InMux I__1765 (
            .O(N__7982),
            .I(N__7976));
    InMux I__1764 (
            .O(N__7981),
            .I(N__7971));
    InMux I__1763 (
            .O(N__7980),
            .I(N__7971));
    InMux I__1762 (
            .O(N__7979),
            .I(N__7968));
    LocalMux I__1761 (
            .O(N__7976),
            .I(N__7961));
    LocalMux I__1760 (
            .O(N__7971),
            .I(N__7961));
    LocalMux I__1759 (
            .O(N__7968),
            .I(N__7961));
    Span4Mux_v I__1758 (
            .O(N__7961),
            .I(N__7957));
    InMux I__1757 (
            .O(N__7960),
            .I(N__7954));
    Odrv4 I__1756 (
            .O(N__7957),
            .I(\Game_Inst.N_16 ));
    LocalMux I__1755 (
            .O(N__7954),
            .I(\Game_Inst.N_16 ));
    IoInMux I__1754 (
            .O(N__7949),
            .I(N__7946));
    LocalMux I__1753 (
            .O(N__7946),
            .I(N__7943));
    IoSpan4Mux I__1752 (
            .O(N__7943),
            .I(N__7940));
    Odrv4 I__1751 (
            .O(N__7940),
            .I(N_87));
    InMux I__1750 (
            .O(N__7937),
            .I(N__7931));
    InMux I__1749 (
            .O(N__7936),
            .I(N__7926));
    InMux I__1748 (
            .O(N__7935),
            .I(N__7926));
    InMux I__1747 (
            .O(N__7934),
            .I(N__7923));
    LocalMux I__1746 (
            .O(N__7931),
            .I(N__7916));
    LocalMux I__1745 (
            .O(N__7926),
            .I(N__7916));
    LocalMux I__1744 (
            .O(N__7923),
            .I(N__7916));
    Odrv4 I__1743 (
            .O(N__7916),
            .I(w_Switch_3));
    InMux I__1742 (
            .O(N__7913),
            .I(N__7910));
    LocalMux I__1741 (
            .O(N__7910),
            .I(N__7907));
    Span4Mux_s3_h I__1740 (
            .O(N__7907),
            .I(N__7904));
    Odrv4 I__1739 (
            .O(N__7904),
            .I(\Debounce_SW3.r_count15_i_a2_0 ));
    CascadeMux I__1738 (
            .O(N__7901),
            .I(N__7898));
    InMux I__1737 (
            .O(N__7898),
            .I(N__7895));
    LocalMux I__1736 (
            .O(N__7895),
            .I(N__7891));
    InMux I__1735 (
            .O(N__7894),
            .I(N__7888));
    Span4Mux_v I__1734 (
            .O(N__7891),
            .I(N__7885));
    LocalMux I__1733 (
            .O(N__7888),
            .I(N__7882));
    Odrv4 I__1732 (
            .O(N__7885),
            .I(i_Switch_3_c));
    Odrv4 I__1731 (
            .O(N__7882),
            .I(i_Switch_3_c));
    InMux I__1730 (
            .O(N__7877),
            .I(N__7874));
    LocalMux I__1729 (
            .O(N__7874),
            .I(N__7871));
    Span4Mux_s3_h I__1728 (
            .O(N__7871),
            .I(N__7868));
    Odrv4 I__1727 (
            .O(N__7868),
            .I(\Debounce_SW3.N_182 ));
    IoInMux I__1726 (
            .O(N__7865),
            .I(N__7862));
    LocalMux I__1725 (
            .O(N__7862),
            .I(\Debounce_SW3.N_40 ));
    InMux I__1724 (
            .O(N__7859),
            .I(N__7856));
    LocalMux I__1723 (
            .O(N__7856),
            .I(\Game_Inst.un1_r_Score_cry_0_THRU_CO ));
    CascadeMux I__1722 (
            .O(N__7853),
            .I(N__7849));
    CascadeMux I__1721 (
            .O(N__7852),
            .I(N__7846));
    InMux I__1720 (
            .O(N__7849),
            .I(N__7832));
    InMux I__1719 (
            .O(N__7846),
            .I(N__7832));
    InMux I__1718 (
            .O(N__7845),
            .I(N__7832));
    InMux I__1717 (
            .O(N__7844),
            .I(N__7832));
    InMux I__1716 (
            .O(N__7843),
            .I(N__7832));
    LocalMux I__1715 (
            .O(N__7832),
            .I(N__7826));
    InMux I__1714 (
            .O(N__7831),
            .I(N__7823));
    InMux I__1713 (
            .O(N__7830),
            .I(N__7820));
    CascadeMux I__1712 (
            .O(N__7829),
            .I(N__7817));
    Span4Mux_s1_v I__1711 (
            .O(N__7826),
            .I(N__7811));
    LocalMux I__1710 (
            .O(N__7823),
            .I(N__7811));
    LocalMux I__1709 (
            .O(N__7820),
            .I(N__7808));
    InMux I__1708 (
            .O(N__7817),
            .I(N__7805));
    CascadeMux I__1707 (
            .O(N__7816),
            .I(N__7802));
    Span4Mux_h I__1706 (
            .O(N__7811),
            .I(N__7798));
    Span4Mux_v I__1705 (
            .O(N__7808),
            .I(N__7793));
    LocalMux I__1704 (
            .O(N__7805),
            .I(N__7793));
    InMux I__1703 (
            .O(N__7802),
            .I(N__7787));
    InMux I__1702 (
            .O(N__7801),
            .I(N__7787));
    Span4Mux_v I__1701 (
            .O(N__7798),
            .I(N__7782));
    Span4Mux_h I__1700 (
            .O(N__7793),
            .I(N__7782));
    InMux I__1699 (
            .O(N__7792),
            .I(N__7779));
    LocalMux I__1698 (
            .O(N__7787),
            .I(w_Score_1));
    Odrv4 I__1697 (
            .O(N__7782),
            .I(w_Score_1));
    LocalMux I__1696 (
            .O(N__7779),
            .I(w_Score_1));
    InMux I__1695 (
            .O(N__7772),
            .I(N__7769));
    LocalMux I__1694 (
            .O(N__7769),
            .I(\Game_Inst.r_Score_RNO_0Z0Z_0 ));
    InMux I__1693 (
            .O(N__7766),
            .I(N__7750));
    InMux I__1692 (
            .O(N__7765),
            .I(N__7750));
    InMux I__1691 (
            .O(N__7764),
            .I(N__7750));
    InMux I__1690 (
            .O(N__7763),
            .I(N__7750));
    InMux I__1689 (
            .O(N__7762),
            .I(N__7750));
    InMux I__1688 (
            .O(N__7761),
            .I(N__7747));
    LocalMux I__1687 (
            .O(N__7750),
            .I(N__7743));
    LocalMux I__1686 (
            .O(N__7747),
            .I(N__7740));
    InMux I__1685 (
            .O(N__7746),
            .I(N__7737));
    Span4Mux_v I__1684 (
            .O(N__7743),
            .I(N__7731));
    Span4Mux_h I__1683 (
            .O(N__7740),
            .I(N__7731));
    LocalMux I__1682 (
            .O(N__7737),
            .I(N__7727));
    InMux I__1681 (
            .O(N__7736),
            .I(N__7724));
    Span4Mux_h I__1680 (
            .O(N__7731),
            .I(N__7720));
    InMux I__1679 (
            .O(N__7730),
            .I(N__7717));
    Span4Mux_v I__1678 (
            .O(N__7727),
            .I(N__7712));
    LocalMux I__1677 (
            .O(N__7724),
            .I(N__7712));
    InMux I__1676 (
            .O(N__7723),
            .I(N__7709));
    Odrv4 I__1675 (
            .O(N__7720),
            .I(w_Score_0));
    LocalMux I__1674 (
            .O(N__7717),
            .I(w_Score_0));
    Odrv4 I__1673 (
            .O(N__7712),
            .I(w_Score_0));
    LocalMux I__1672 (
            .O(N__7709),
            .I(w_Score_0));
    InMux I__1671 (
            .O(N__7700),
            .I(N__7693));
    InMux I__1670 (
            .O(N__7699),
            .I(N__7690));
    InMux I__1669 (
            .O(N__7698),
            .I(N__7687));
    InMux I__1668 (
            .O(N__7697),
            .I(N__7681));
    InMux I__1667 (
            .O(N__7696),
            .I(N__7681));
    LocalMux I__1666 (
            .O(N__7693),
            .I(N__7676));
    LocalMux I__1665 (
            .O(N__7690),
            .I(N__7671));
    LocalMux I__1664 (
            .O(N__7687),
            .I(N__7671));
    InMux I__1663 (
            .O(N__7686),
            .I(N__7668));
    LocalMux I__1662 (
            .O(N__7681),
            .I(N__7665));
    InMux I__1661 (
            .O(N__7680),
            .I(N__7660));
    InMux I__1660 (
            .O(N__7679),
            .I(N__7660));
    Span4Mux_v I__1659 (
            .O(N__7676),
            .I(N__7645));
    Span4Mux_v I__1658 (
            .O(N__7671),
            .I(N__7645));
    LocalMux I__1657 (
            .O(N__7668),
            .I(N__7645));
    Span4Mux_v I__1656 (
            .O(N__7665),
            .I(N__7642));
    LocalMux I__1655 (
            .O(N__7660),
            .I(N__7639));
    InMux I__1654 (
            .O(N__7659),
            .I(N__7632));
    InMux I__1653 (
            .O(N__7658),
            .I(N__7632));
    InMux I__1652 (
            .O(N__7657),
            .I(N__7632));
    InMux I__1651 (
            .O(N__7656),
            .I(N__7625));
    InMux I__1650 (
            .O(N__7655),
            .I(N__7625));
    InMux I__1649 (
            .O(N__7654),
            .I(N__7625));
    InMux I__1648 (
            .O(N__7653),
            .I(N__7620));
    InMux I__1647 (
            .O(N__7652),
            .I(N__7620));
    Span4Mux_h I__1646 (
            .O(N__7645),
            .I(N__7617));
    Odrv4 I__1645 (
            .O(N__7642),
            .I(\Game_Inst.r_SM_MainZ0Z_0 ));
    Odrv4 I__1644 (
            .O(N__7639),
            .I(\Game_Inst.r_SM_MainZ0Z_0 ));
    LocalMux I__1643 (
            .O(N__7632),
            .I(\Game_Inst.r_SM_MainZ0Z_0 ));
    LocalMux I__1642 (
            .O(N__7625),
            .I(\Game_Inst.r_SM_MainZ0Z_0 ));
    LocalMux I__1641 (
            .O(N__7620),
            .I(\Game_Inst.r_SM_MainZ0Z_0 ));
    Odrv4 I__1640 (
            .O(N__7617),
            .I(\Game_Inst.r_SM_MainZ0Z_0 ));
    InMux I__1639 (
            .O(N__7604),
            .I(N__7596));
    InMux I__1638 (
            .O(N__7603),
            .I(N__7590));
    InMux I__1637 (
            .O(N__7602),
            .I(N__7587));
    InMux I__1636 (
            .O(N__7601),
            .I(N__7584));
    InMux I__1635 (
            .O(N__7600),
            .I(N__7580));
    InMux I__1634 (
            .O(N__7599),
            .I(N__7577));
    LocalMux I__1633 (
            .O(N__7596),
            .I(N__7573));
    InMux I__1632 (
            .O(N__7595),
            .I(N__7568));
    InMux I__1631 (
            .O(N__7594),
            .I(N__7568));
    CascadeMux I__1630 (
            .O(N__7593),
            .I(N__7563));
    LocalMux I__1629 (
            .O(N__7590),
            .I(N__7560));
    LocalMux I__1628 (
            .O(N__7587),
            .I(N__7555));
    LocalMux I__1627 (
            .O(N__7584),
            .I(N__7552));
    CascadeMux I__1626 (
            .O(N__7583),
            .I(N__7549));
    LocalMux I__1625 (
            .O(N__7580),
            .I(N__7544));
    LocalMux I__1624 (
            .O(N__7577),
            .I(N__7544));
    CascadeMux I__1623 (
            .O(N__7576),
            .I(N__7541));
    Span4Mux_v I__1622 (
            .O(N__7573),
            .I(N__7535));
    LocalMux I__1621 (
            .O(N__7568),
            .I(N__7535));
    InMux I__1620 (
            .O(N__7567),
            .I(N__7528));
    InMux I__1619 (
            .O(N__7566),
            .I(N__7528));
    InMux I__1618 (
            .O(N__7563),
            .I(N__7528));
    Span4Mux_h I__1617 (
            .O(N__7560),
            .I(N__7525));
    InMux I__1616 (
            .O(N__7559),
            .I(N__7522));
    InMux I__1615 (
            .O(N__7558),
            .I(N__7519));
    Span4Mux_v I__1614 (
            .O(N__7555),
            .I(N__7514));
    Span4Mux_h I__1613 (
            .O(N__7552),
            .I(N__7514));
    InMux I__1612 (
            .O(N__7549),
            .I(N__7511));
    Span4Mux_h I__1611 (
            .O(N__7544),
            .I(N__7508));
    InMux I__1610 (
            .O(N__7541),
            .I(N__7503));
    InMux I__1609 (
            .O(N__7540),
            .I(N__7503));
    Odrv4 I__1608 (
            .O(N__7535),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    LocalMux I__1607 (
            .O(N__7528),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    Odrv4 I__1606 (
            .O(N__7525),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    LocalMux I__1605 (
            .O(N__7522),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    LocalMux I__1604 (
            .O(N__7519),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    Odrv4 I__1603 (
            .O(N__7514),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    LocalMux I__1602 (
            .O(N__7511),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    Odrv4 I__1601 (
            .O(N__7508),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    LocalMux I__1600 (
            .O(N__7503),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    InMux I__1599 (
            .O(N__7484),
            .I(N__7480));
    InMux I__1598 (
            .O(N__7483),
            .I(N__7476));
    LocalMux I__1597 (
            .O(N__7480),
            .I(N__7472));
    InMux I__1596 (
            .O(N__7479),
            .I(N__7469));
    LocalMux I__1595 (
            .O(N__7476),
            .I(N__7464));
    CascadeMux I__1594 (
            .O(N__7475),
            .I(N__7461));
    Span4Mux_v I__1593 (
            .O(N__7472),
            .I(N__7455));
    LocalMux I__1592 (
            .O(N__7469),
            .I(N__7455));
    InMux I__1591 (
            .O(N__7468),
            .I(N__7452));
    InMux I__1590 (
            .O(N__7467),
            .I(N__7449));
    Span4Mux_v I__1589 (
            .O(N__7464),
            .I(N__7446));
    InMux I__1588 (
            .O(N__7461),
            .I(N__7443));
    InMux I__1587 (
            .O(N__7460),
            .I(N__7440));
    Span4Mux_v I__1586 (
            .O(N__7455),
            .I(N__7437));
    LocalMux I__1585 (
            .O(N__7452),
            .I(N__7434));
    LocalMux I__1584 (
            .O(N__7449),
            .I(N__7431));
    Odrv4 I__1583 (
            .O(N__7446),
            .I(\Game_Inst.N_291 ));
    LocalMux I__1582 (
            .O(N__7443),
            .I(\Game_Inst.N_291 ));
    LocalMux I__1581 (
            .O(N__7440),
            .I(\Game_Inst.N_291 ));
    Odrv4 I__1580 (
            .O(N__7437),
            .I(\Game_Inst.N_291 ));
    Odrv4 I__1579 (
            .O(N__7434),
            .I(\Game_Inst.N_291 ));
    Odrv12 I__1578 (
            .O(N__7431),
            .I(\Game_Inst.N_291 ));
    InMux I__1577 (
            .O(N__7418),
            .I(N__7410));
    InMux I__1576 (
            .O(N__7417),
            .I(N__7407));
    CascadeMux I__1575 (
            .O(N__7416),
            .I(N__7399));
    CascadeMux I__1574 (
            .O(N__7415),
            .I(N__7394));
    InMux I__1573 (
            .O(N__7414),
            .I(N__7388));
    InMux I__1572 (
            .O(N__7413),
            .I(N__7388));
    LocalMux I__1571 (
            .O(N__7410),
            .I(N__7381));
    LocalMux I__1570 (
            .O(N__7407),
            .I(N__7381));
    InMux I__1569 (
            .O(N__7406),
            .I(N__7376));
    InMux I__1568 (
            .O(N__7405),
            .I(N__7376));
    InMux I__1567 (
            .O(N__7404),
            .I(N__7369));
    InMux I__1566 (
            .O(N__7403),
            .I(N__7369));
    InMux I__1565 (
            .O(N__7402),
            .I(N__7369));
    InMux I__1564 (
            .O(N__7399),
            .I(N__7364));
    InMux I__1563 (
            .O(N__7398),
            .I(N__7364));
    InMux I__1562 (
            .O(N__7397),
            .I(N__7361));
    InMux I__1561 (
            .O(N__7394),
            .I(N__7356));
    InMux I__1560 (
            .O(N__7393),
            .I(N__7356));
    LocalMux I__1559 (
            .O(N__7388),
            .I(N__7353));
    InMux I__1558 (
            .O(N__7387),
            .I(N__7348));
    InMux I__1557 (
            .O(N__7386),
            .I(N__7348));
    Span4Mux_h I__1556 (
            .O(N__7381),
            .I(N__7343));
    LocalMux I__1555 (
            .O(N__7376),
            .I(N__7343));
    LocalMux I__1554 (
            .O(N__7369),
            .I(N__7340));
    LocalMux I__1553 (
            .O(N__7364),
            .I(N__7337));
    LocalMux I__1552 (
            .O(N__7361),
            .I(\Game_Inst.r_SM_MainZ0Z_1 ));
    LocalMux I__1551 (
            .O(N__7356),
            .I(\Game_Inst.r_SM_MainZ0Z_1 ));
    Odrv4 I__1550 (
            .O(N__7353),
            .I(\Game_Inst.r_SM_MainZ0Z_1 ));
    LocalMux I__1549 (
            .O(N__7348),
            .I(\Game_Inst.r_SM_MainZ0Z_1 ));
    Odrv4 I__1548 (
            .O(N__7343),
            .I(\Game_Inst.r_SM_MainZ0Z_1 ));
    Odrv12 I__1547 (
            .O(N__7340),
            .I(\Game_Inst.r_SM_MainZ0Z_1 ));
    Odrv4 I__1546 (
            .O(N__7337),
            .I(\Game_Inst.r_SM_MainZ0Z_1 ));
    InMux I__1545 (
            .O(N__7322),
            .I(N__7319));
    LocalMux I__1544 (
            .O(N__7319),
            .I(\Game_Inst.N_241 ));
    InMux I__1543 (
            .O(N__7316),
            .I(N__7310));
    InMux I__1542 (
            .O(N__7315),
            .I(N__7303));
    InMux I__1541 (
            .O(N__7314),
            .I(N__7303));
    InMux I__1540 (
            .O(N__7313),
            .I(N__7303));
    LocalMux I__1539 (
            .O(N__7310),
            .I(N__7300));
    LocalMux I__1538 (
            .O(N__7303),
            .I(N__7296));
    Span4Mux_h I__1537 (
            .O(N__7300),
            .I(N__7293));
    InMux I__1536 (
            .O(N__7299),
            .I(N__7290));
    Odrv4 I__1535 (
            .O(N__7296),
            .I(\Game_Inst.r_Score_0_sqmuxa ));
    Odrv4 I__1534 (
            .O(N__7293),
            .I(\Game_Inst.r_Score_0_sqmuxa ));
    LocalMux I__1533 (
            .O(N__7290),
            .I(\Game_Inst.r_Score_0_sqmuxa ));
    CascadeMux I__1532 (
            .O(N__7283),
            .I(N__7278));
    InMux I__1531 (
            .O(N__7282),
            .I(N__7270));
    InMux I__1530 (
            .O(N__7281),
            .I(N__7270));
    InMux I__1529 (
            .O(N__7278),
            .I(N__7270));
    InMux I__1528 (
            .O(N__7277),
            .I(N__7267));
    LocalMux I__1527 (
            .O(N__7270),
            .I(\Game_Inst.un1_r_SM_Main_0 ));
    LocalMux I__1526 (
            .O(N__7267),
            .I(\Game_Inst.un1_r_SM_Main_0 ));
    CascadeMux I__1525 (
            .O(N__7262),
            .I(\Game_Inst.N_241_cascade_ ));
    InMux I__1524 (
            .O(N__7259),
            .I(N__7256));
    LocalMux I__1523 (
            .O(N__7256),
            .I(\Game_Inst.r_Score_RNO_0Z0Z_2 ));
    InMux I__1522 (
            .O(N__7253),
            .I(N__7238));
    InMux I__1521 (
            .O(N__7252),
            .I(N__7238));
    InMux I__1520 (
            .O(N__7251),
            .I(N__7238));
    InMux I__1519 (
            .O(N__7250),
            .I(N__7238));
    InMux I__1518 (
            .O(N__7249),
            .I(N__7238));
    LocalMux I__1517 (
            .O(N__7238),
            .I(N__7231));
    InMux I__1516 (
            .O(N__7237),
            .I(N__7228));
    InMux I__1515 (
            .O(N__7236),
            .I(N__7225));
    InMux I__1514 (
            .O(N__7235),
            .I(N__7222));
    CascadeMux I__1513 (
            .O(N__7234),
            .I(N__7219));
    Span4Mux_s1_v I__1512 (
            .O(N__7231),
            .I(N__7214));
    LocalMux I__1511 (
            .O(N__7228),
            .I(N__7214));
    LocalMux I__1510 (
            .O(N__7225),
            .I(N__7211));
    LocalMux I__1509 (
            .O(N__7222),
            .I(N__7207));
    InMux I__1508 (
            .O(N__7219),
            .I(N__7204));
    Span4Mux_h I__1507 (
            .O(N__7214),
            .I(N__7199));
    Span4Mux_h I__1506 (
            .O(N__7211),
            .I(N__7199));
    InMux I__1505 (
            .O(N__7210),
            .I(N__7196));
    Odrv12 I__1504 (
            .O(N__7207),
            .I(w_Score_2));
    LocalMux I__1503 (
            .O(N__7204),
            .I(w_Score_2));
    Odrv4 I__1502 (
            .O(N__7199),
            .I(w_Score_2));
    LocalMux I__1501 (
            .O(N__7196),
            .I(w_Score_2));
    InMux I__1500 (
            .O(N__7187),
            .I(N__7183));
    InMux I__1499 (
            .O(N__7186),
            .I(N__7180));
    LocalMux I__1498 (
            .O(N__7183),
            .I(\Game_Inst.w_LFSR_Data_8 ));
    LocalMux I__1497 (
            .O(N__7180),
            .I(\Game_Inst.w_LFSR_Data_8 ));
    InMux I__1496 (
            .O(N__7175),
            .I(N__7171));
    InMux I__1495 (
            .O(N__7174),
            .I(N__7168));
    LocalMux I__1494 (
            .O(N__7171),
            .I(N__7165));
    LocalMux I__1493 (
            .O(N__7168),
            .I(\Game_Inst.w_LFSR_Data_9 ));
    Odrv4 I__1492 (
            .O(N__7165),
            .I(\Game_Inst.w_LFSR_Data_9 ));
    InMux I__1491 (
            .O(N__7160),
            .I(N__7157));
    LocalMux I__1490 (
            .O(N__7157),
            .I(N__7153));
    InMux I__1489 (
            .O(N__7156),
            .I(N__7150));
    Span4Mux_h I__1488 (
            .O(N__7153),
            .I(N__7145));
    LocalMux I__1487 (
            .O(N__7150),
            .I(N__7145));
    Sp12to4 I__1486 (
            .O(N__7145),
            .I(N__7142));
    Span12Mux_v I__1485 (
            .O(N__7142),
            .I(N__7139));
    Odrv12 I__1484 (
            .O(N__7139),
            .I(i_Switch_2_c));
    CEMux I__1483 (
            .O(N__7136),
            .I(N__7133));
    LocalMux I__1482 (
            .O(N__7133),
            .I(N__7130));
    Odrv12 I__1481 (
            .O(N__7130),
            .I(\Debounce_SW2.r_State_e_0_RNOZ0Z_0 ));
    CEMux I__1480 (
            .O(N__7127),
            .I(N__7124));
    LocalMux I__1479 (
            .O(N__7124),
            .I(N__7121));
    Span4Mux_s3_h I__1478 (
            .O(N__7121),
            .I(N__7118));
    Odrv4 I__1477 (
            .O(N__7118),
            .I(\Debounce_SW3.r_State_e_0_RNO_1 ));
    CascadeMux I__1476 (
            .O(N__7115),
            .I(N__7109));
    InMux I__1475 (
            .O(N__7114),
            .I(N__7106));
    InMux I__1474 (
            .O(N__7113),
            .I(N__7102));
    InMux I__1473 (
            .O(N__7112),
            .I(N__7099));
    InMux I__1472 (
            .O(N__7109),
            .I(N__7095));
    LocalMux I__1471 (
            .O(N__7106),
            .I(N__7090));
    InMux I__1470 (
            .O(N__7105),
            .I(N__7087));
    LocalMux I__1469 (
            .O(N__7102),
            .I(N__7082));
    LocalMux I__1468 (
            .O(N__7099),
            .I(N__7082));
    InMux I__1467 (
            .O(N__7098),
            .I(N__7079));
    LocalMux I__1466 (
            .O(N__7095),
            .I(N__7076));
    InMux I__1465 (
            .O(N__7094),
            .I(N__7071));
    InMux I__1464 (
            .O(N__7093),
            .I(N__7071));
    Span4Mux_v I__1463 (
            .O(N__7090),
            .I(N__7066));
    LocalMux I__1462 (
            .O(N__7087),
            .I(N__7066));
    Span4Mux_h I__1461 (
            .O(N__7082),
            .I(N__7061));
    LocalMux I__1460 (
            .O(N__7079),
            .I(N__7061));
    Odrv12 I__1459 (
            .O(N__7076),
            .I(w_Switch_1));
    LocalMux I__1458 (
            .O(N__7071),
            .I(w_Switch_1));
    Odrv4 I__1457 (
            .O(N__7066),
            .I(w_Switch_1));
    Odrv4 I__1456 (
            .O(N__7061),
            .I(w_Switch_1));
    IoInMux I__1455 (
            .O(N__7052),
            .I(N__7049));
    LocalMux I__1454 (
            .O(N__7049),
            .I(N__7046));
    IoSpan4Mux I__1453 (
            .O(N__7046),
            .I(N__7043));
    Odrv4 I__1452 (
            .O(N__7043),
            .I(N_70));
    InMux I__1451 (
            .O(N__7040),
            .I(N__7036));
    InMux I__1450 (
            .O(N__7039),
            .I(N__7033));
    LocalMux I__1449 (
            .O(N__7036),
            .I(\Game_Inst.w_LFSR_Data_11 ));
    LocalMux I__1448 (
            .O(N__7033),
            .I(\Game_Inst.w_LFSR_Data_11 ));
    InMux I__1447 (
            .O(N__7028),
            .I(N__7025));
    LocalMux I__1446 (
            .O(N__7025),
            .I(N__7022));
    Span4Mux_v I__1445 (
            .O(N__7022),
            .I(N__7018));
    InMux I__1444 (
            .O(N__7021),
            .I(N__7015));
    Odrv4 I__1443 (
            .O(N__7018),
            .I(\Game_Inst.w_LFSR_Data_12 ));
    LocalMux I__1442 (
            .O(N__7015),
            .I(\Game_Inst.w_LFSR_Data_12 ));
    InMux I__1441 (
            .O(N__7010),
            .I(N__7007));
    LocalMux I__1440 (
            .O(N__7007),
            .I(N__7004));
    Span4Mux_v I__1439 (
            .O(N__7004),
            .I(N__7000));
    InMux I__1438 (
            .O(N__7003),
            .I(N__6997));
    Odrv4 I__1437 (
            .O(N__7000),
            .I(\Game_Inst.w_LFSR_Data_13 ));
    LocalMux I__1436 (
            .O(N__6997),
            .I(\Game_Inst.w_LFSR_Data_13 ));
    InMux I__1435 (
            .O(N__6992),
            .I(N__6988));
    InMux I__1434 (
            .O(N__6991),
            .I(N__6985));
    LocalMux I__1433 (
            .O(N__6988),
            .I(\Game_Inst.w_LFSR_Data_10 ));
    LocalMux I__1432 (
            .O(N__6985),
            .I(\Game_Inst.w_LFSR_Data_10 ));
    InMux I__1431 (
            .O(N__6980),
            .I(\Game_Inst.un1_r_Score_cry_0 ));
    InMux I__1430 (
            .O(N__6977),
            .I(\Game_Inst.un1_r_Score_cry_1 ));
    InMux I__1429 (
            .O(N__6974),
            .I(\Game_Inst.un1_r_Score_cry_2 ));
    CascadeMux I__1428 (
            .O(N__6971),
            .I(N__6964));
    CascadeMux I__1427 (
            .O(N__6970),
            .I(N__6961));
    CascadeMux I__1426 (
            .O(N__6969),
            .I(N__6958));
    InMux I__1425 (
            .O(N__6968),
            .I(N__6945));
    InMux I__1424 (
            .O(N__6967),
            .I(N__6945));
    InMux I__1423 (
            .O(N__6964),
            .I(N__6945));
    InMux I__1422 (
            .O(N__6961),
            .I(N__6945));
    InMux I__1421 (
            .O(N__6958),
            .I(N__6945));
    CascadeMux I__1420 (
            .O(N__6957),
            .I(N__6942));
    CascadeMux I__1419 (
            .O(N__6956),
            .I(N__6939));
    LocalMux I__1418 (
            .O(N__6945),
            .I(N__6935));
    InMux I__1417 (
            .O(N__6942),
            .I(N__6932));
    InMux I__1416 (
            .O(N__6939),
            .I(N__6929));
    CascadeMux I__1415 (
            .O(N__6938),
            .I(N__6925));
    Span4Mux_s1_v I__1414 (
            .O(N__6935),
            .I(N__6920));
    LocalMux I__1413 (
            .O(N__6932),
            .I(N__6920));
    LocalMux I__1412 (
            .O(N__6929),
            .I(N__6917));
    InMux I__1411 (
            .O(N__6928),
            .I(N__6914));
    InMux I__1410 (
            .O(N__6925),
            .I(N__6910));
    Span4Mux_h I__1409 (
            .O(N__6920),
            .I(N__6907));
    Span4Mux_v I__1408 (
            .O(N__6917),
            .I(N__6902));
    LocalMux I__1407 (
            .O(N__6914),
            .I(N__6902));
    CascadeMux I__1406 (
            .O(N__6913),
            .I(N__6899));
    LocalMux I__1405 (
            .O(N__6910),
            .I(N__6892));
    Span4Mux_v I__1404 (
            .O(N__6907),
            .I(N__6892));
    Span4Mux_h I__1403 (
            .O(N__6902),
            .I(N__6892));
    InMux I__1402 (
            .O(N__6899),
            .I(N__6889));
    Odrv4 I__1401 (
            .O(N__6892),
            .I(w_Score_3));
    LocalMux I__1400 (
            .O(N__6889),
            .I(w_Score_3));
    CascadeMux I__1399 (
            .O(N__6884),
            .I(\Game_Inst.N_291_cascade_ ));
    CascadeMux I__1398 (
            .O(N__6881),
            .I(N__6877));
    InMux I__1397 (
            .O(N__6880),
            .I(N__6874));
    InMux I__1396 (
            .O(N__6877),
            .I(N__6871));
    LocalMux I__1395 (
            .O(N__6874),
            .I(\Game_Inst.N_68_i ));
    LocalMux I__1394 (
            .O(N__6871),
            .I(\Game_Inst.N_68_i ));
    CascadeMux I__1393 (
            .O(N__6866),
            .I(N__6861));
    InMux I__1392 (
            .O(N__6865),
            .I(N__6858));
    InMux I__1391 (
            .O(N__6864),
            .I(N__6855));
    InMux I__1390 (
            .O(N__6861),
            .I(N__6852));
    LocalMux I__1389 (
            .O(N__6858),
            .I(\Debounce_SW3.r_CountZ0Z_13 ));
    LocalMux I__1388 (
            .O(N__6855),
            .I(\Debounce_SW3.r_CountZ0Z_13 ));
    LocalMux I__1387 (
            .O(N__6852),
            .I(\Debounce_SW3.r_CountZ0Z_13 ));
    InMux I__1386 (
            .O(N__6845),
            .I(\Debounce_SW3.un2_r_count_cry_12 ));
    InMux I__1385 (
            .O(N__6842),
            .I(N__6838));
    InMux I__1384 (
            .O(N__6841),
            .I(N__6835));
    LocalMux I__1383 (
            .O(N__6838),
            .I(\Debounce_SW3.r_CountZ0Z_14 ));
    LocalMux I__1382 (
            .O(N__6835),
            .I(\Debounce_SW3.r_CountZ0Z_14 ));
    InMux I__1381 (
            .O(N__6830),
            .I(\Debounce_SW3.un2_r_count_cry_13 ));
    InMux I__1380 (
            .O(N__6827),
            .I(N__6823));
    InMux I__1379 (
            .O(N__6826),
            .I(N__6820));
    LocalMux I__1378 (
            .O(N__6823),
            .I(\Debounce_SW3.r_CountZ0Z_15 ));
    LocalMux I__1377 (
            .O(N__6820),
            .I(\Debounce_SW3.r_CountZ0Z_15 ));
    InMux I__1376 (
            .O(N__6815),
            .I(\Debounce_SW3.un2_r_count_cry_14 ));
    InMux I__1375 (
            .O(N__6812),
            .I(N__6808));
    InMux I__1374 (
            .O(N__6811),
            .I(N__6805));
    LocalMux I__1373 (
            .O(N__6808),
            .I(\Debounce_SW3.r_CountZ0Z_16 ));
    LocalMux I__1372 (
            .O(N__6805),
            .I(\Debounce_SW3.r_CountZ0Z_16 ));
    InMux I__1371 (
            .O(N__6800),
            .I(\Debounce_SW3.un2_r_count_cry_15 ));
    InMux I__1370 (
            .O(N__6797),
            .I(bfn_9_7_0_));
    CascadeMux I__1369 (
            .O(N__6794),
            .I(N__6791));
    InMux I__1368 (
            .O(N__6791),
            .I(N__6787));
    InMux I__1367 (
            .O(N__6790),
            .I(N__6784));
    LocalMux I__1366 (
            .O(N__6787),
            .I(N__6781));
    LocalMux I__1365 (
            .O(N__6784),
            .I(\Debounce_SW3.r_CountZ0Z_17 ));
    Odrv4 I__1364 (
            .O(N__6781),
            .I(\Debounce_SW3.r_CountZ0Z_17 ));
    SRMux I__1363 (
            .O(N__6776),
            .I(N__6764));
    SRMux I__1362 (
            .O(N__6775),
            .I(N__6764));
    SRMux I__1361 (
            .O(N__6774),
            .I(N__6764));
    SRMux I__1360 (
            .O(N__6773),
            .I(N__6764));
    GlobalMux I__1359 (
            .O(N__6764),
            .I(N__6761));
    gio2CtrlBuf I__1358 (
            .O(N__6761),
            .I(\Debounce_SW3.N_40_g ));
    InMux I__1357 (
            .O(N__6758),
            .I(N__6755));
    LocalMux I__1356 (
            .O(N__6755),
            .I(N__6751));
    InMux I__1355 (
            .O(N__6754),
            .I(N__6748));
    Span4Mux_h I__1354 (
            .O(N__6751),
            .I(N__6743));
    LocalMux I__1353 (
            .O(N__6748),
            .I(N__6743));
    Span4Mux_v I__1352 (
            .O(N__6743),
            .I(N__6740));
    Odrv4 I__1351 (
            .O(N__6740),
            .I(i_Switch_1_c));
    CEMux I__1350 (
            .O(N__6737),
            .I(N__6734));
    LocalMux I__1349 (
            .O(N__6734),
            .I(N__6731));
    Odrv4 I__1348 (
            .O(N__6731),
            .I(\Debounce_SW1.r_State_e_0_RNOZ0 ));
    InMux I__1347 (
            .O(N__6728),
            .I(N__6724));
    InMux I__1346 (
            .O(N__6727),
            .I(N__6721));
    LocalMux I__1345 (
            .O(N__6724),
            .I(\Debounce_SW3.r_CountZ0Z_4 ));
    LocalMux I__1344 (
            .O(N__6721),
            .I(\Debounce_SW3.r_CountZ0Z_4 ));
    InMux I__1343 (
            .O(N__6716),
            .I(\Debounce_SW3.un2_r_count_cry_3 ));
    InMux I__1342 (
            .O(N__6713),
            .I(N__6709));
    InMux I__1341 (
            .O(N__6712),
            .I(N__6706));
    LocalMux I__1340 (
            .O(N__6709),
            .I(\Debounce_SW3.r_CountZ0Z_5 ));
    LocalMux I__1339 (
            .O(N__6706),
            .I(\Debounce_SW3.r_CountZ0Z_5 ));
    InMux I__1338 (
            .O(N__6701),
            .I(\Debounce_SW3.un2_r_count_cry_4 ));
    InMux I__1337 (
            .O(N__6698),
            .I(N__6694));
    InMux I__1336 (
            .O(N__6697),
            .I(N__6691));
    LocalMux I__1335 (
            .O(N__6694),
            .I(\Debounce_SW3.r_CountZ0Z_6 ));
    LocalMux I__1334 (
            .O(N__6691),
            .I(\Debounce_SW3.r_CountZ0Z_6 ));
    InMux I__1333 (
            .O(N__6686),
            .I(\Debounce_SW3.un2_r_count_cry_5 ));
    InMux I__1332 (
            .O(N__6683),
            .I(N__6678));
    InMux I__1331 (
            .O(N__6682),
            .I(N__6673));
    InMux I__1330 (
            .O(N__6681),
            .I(N__6673));
    LocalMux I__1329 (
            .O(N__6678),
            .I(\Debounce_SW3.r_CountZ0Z_7 ));
    LocalMux I__1328 (
            .O(N__6673),
            .I(\Debounce_SW3.r_CountZ0Z_7 ));
    InMux I__1327 (
            .O(N__6668),
            .I(\Debounce_SW3.un2_r_count_cry_6 ));
    InMux I__1326 (
            .O(N__6665),
            .I(N__6661));
    InMux I__1325 (
            .O(N__6664),
            .I(N__6658));
    LocalMux I__1324 (
            .O(N__6661),
            .I(\Debounce_SW3.r_CountZ0Z_8 ));
    LocalMux I__1323 (
            .O(N__6658),
            .I(\Debounce_SW3.r_CountZ0Z_8 ));
    InMux I__1322 (
            .O(N__6653),
            .I(\Debounce_SW3.un2_r_count_cry_7 ));
    InMux I__1321 (
            .O(N__6650),
            .I(N__6646));
    InMux I__1320 (
            .O(N__6649),
            .I(N__6643));
    LocalMux I__1319 (
            .O(N__6646),
            .I(\Debounce_SW3.r_CountZ0Z_9 ));
    LocalMux I__1318 (
            .O(N__6643),
            .I(\Debounce_SW3.r_CountZ0Z_9 ));
    InMux I__1317 (
            .O(N__6638),
            .I(bfn_9_6_0_));
    InMux I__1316 (
            .O(N__6635),
            .I(N__6631));
    InMux I__1315 (
            .O(N__6634),
            .I(N__6628));
    LocalMux I__1314 (
            .O(N__6631),
            .I(N__6625));
    LocalMux I__1313 (
            .O(N__6628),
            .I(\Debounce_SW3.r_CountZ0Z_10 ));
    Odrv4 I__1312 (
            .O(N__6625),
            .I(\Debounce_SW3.r_CountZ0Z_10 ));
    InMux I__1311 (
            .O(N__6620),
            .I(\Debounce_SW3.un2_r_count_cry_9 ));
    CascadeMux I__1310 (
            .O(N__6617),
            .I(N__6613));
    InMux I__1309 (
            .O(N__6616),
            .I(N__6610));
    InMux I__1308 (
            .O(N__6613),
            .I(N__6607));
    LocalMux I__1307 (
            .O(N__6610),
            .I(\Debounce_SW3.r_CountZ0Z_11 ));
    LocalMux I__1306 (
            .O(N__6607),
            .I(\Debounce_SW3.r_CountZ0Z_11 ));
    InMux I__1305 (
            .O(N__6602),
            .I(\Debounce_SW3.un2_r_count_cry_10 ));
    InMux I__1304 (
            .O(N__6599),
            .I(N__6594));
    InMux I__1303 (
            .O(N__6598),
            .I(N__6589));
    InMux I__1302 (
            .O(N__6597),
            .I(N__6589));
    LocalMux I__1301 (
            .O(N__6594),
            .I(\Debounce_SW3.r_CountZ0Z_12 ));
    LocalMux I__1300 (
            .O(N__6589),
            .I(\Debounce_SW3.r_CountZ0Z_12 ));
    InMux I__1299 (
            .O(N__6584),
            .I(\Debounce_SW3.un2_r_count_cry_11 ));
    InMux I__1298 (
            .O(N__6581),
            .I(N__6576));
    InMux I__1297 (
            .O(N__6580),
            .I(N__6571));
    InMux I__1296 (
            .O(N__6579),
            .I(N__6571));
    LocalMux I__1295 (
            .O(N__6576),
            .I(\Debounce_SW2.r_CountZ0Z_7 ));
    LocalMux I__1294 (
            .O(N__6571),
            .I(\Debounce_SW2.r_CountZ0Z_7 ));
    CascadeMux I__1293 (
            .O(N__6566),
            .I(\Debounce_SW2.N_147_cascade_ ));
    InMux I__1292 (
            .O(N__6563),
            .I(N__6560));
    LocalMux I__1291 (
            .O(N__6560),
            .I(\Debounce_SW2.N_286 ));
    InMux I__1290 (
            .O(N__6557),
            .I(N__6553));
    InMux I__1289 (
            .O(N__6556),
            .I(N__6550));
    LocalMux I__1288 (
            .O(N__6553),
            .I(\Debounce_SW2.r_CountZ0Z_2 ));
    LocalMux I__1287 (
            .O(N__6550),
            .I(\Debounce_SW2.r_CountZ0Z_2 ));
    CascadeMux I__1286 (
            .O(N__6545),
            .I(N__6541));
    InMux I__1285 (
            .O(N__6544),
            .I(N__6538));
    InMux I__1284 (
            .O(N__6541),
            .I(N__6535));
    LocalMux I__1283 (
            .O(N__6538),
            .I(\Debounce_SW2.r_CountZ0Z_3 ));
    LocalMux I__1282 (
            .O(N__6535),
            .I(\Debounce_SW2.r_CountZ0Z_3 ));
    InMux I__1281 (
            .O(N__6530),
            .I(N__6524));
    InMux I__1280 (
            .O(N__6529),
            .I(N__6524));
    LocalMux I__1279 (
            .O(N__6524),
            .I(\Debounce_SW2.un9_r_count_10 ));
    InMux I__1278 (
            .O(N__6521),
            .I(N__6517));
    InMux I__1277 (
            .O(N__6520),
            .I(N__6514));
    LocalMux I__1276 (
            .O(N__6517),
            .I(\Debounce_SW2.r_CountZ0Z_16 ));
    LocalMux I__1275 (
            .O(N__6514),
            .I(\Debounce_SW2.r_CountZ0Z_16 ));
    InMux I__1274 (
            .O(N__6509),
            .I(N__6505));
    InMux I__1273 (
            .O(N__6508),
            .I(N__6502));
    LocalMux I__1272 (
            .O(N__6505),
            .I(\Debounce_SW2.r_CountZ0Z_15 ));
    LocalMux I__1271 (
            .O(N__6502),
            .I(\Debounce_SW2.r_CountZ0Z_15 ));
    CascadeMux I__1270 (
            .O(N__6497),
            .I(N__6493));
    InMux I__1269 (
            .O(N__6496),
            .I(N__6490));
    InMux I__1268 (
            .O(N__6493),
            .I(N__6487));
    LocalMux I__1267 (
            .O(N__6490),
            .I(\Debounce_SW2.r_CountZ0Z_17 ));
    LocalMux I__1266 (
            .O(N__6487),
            .I(\Debounce_SW2.r_CountZ0Z_17 ));
    InMux I__1265 (
            .O(N__6482),
            .I(N__6478));
    InMux I__1264 (
            .O(N__6481),
            .I(N__6475));
    LocalMux I__1263 (
            .O(N__6478),
            .I(\Debounce_SW2.r_CountZ0Z_14 ));
    LocalMux I__1262 (
            .O(N__6475),
            .I(\Debounce_SW2.r_CountZ0Z_14 ));
    InMux I__1261 (
            .O(N__6470),
            .I(N__6464));
    InMux I__1260 (
            .O(N__6469),
            .I(N__6464));
    LocalMux I__1259 (
            .O(N__6464),
            .I(\Debounce_SW2.r_count15_i_a2_0 ));
    CascadeMux I__1258 (
            .O(N__6461),
            .I(N__6458));
    InMux I__1257 (
            .O(N__6458),
            .I(N__6454));
    InMux I__1256 (
            .O(N__6457),
            .I(N__6450));
    LocalMux I__1255 (
            .O(N__6454),
            .I(N__6447));
    InMux I__1254 (
            .O(N__6453),
            .I(N__6444));
    LocalMux I__1253 (
            .O(N__6450),
            .I(\Debounce_SW2.r_CountZ0Z_1 ));
    Odrv4 I__1252 (
            .O(N__6447),
            .I(\Debounce_SW2.r_CountZ0Z_1 ));
    LocalMux I__1251 (
            .O(N__6444),
            .I(\Debounce_SW2.r_CountZ0Z_1 ));
    InMux I__1250 (
            .O(N__6437),
            .I(N__6432));
    InMux I__1249 (
            .O(N__6436),
            .I(N__6426));
    InMux I__1248 (
            .O(N__6435),
            .I(N__6426));
    LocalMux I__1247 (
            .O(N__6432),
            .I(N__6423));
    InMux I__1246 (
            .O(N__6431),
            .I(N__6420));
    LocalMux I__1245 (
            .O(N__6426),
            .I(\Debounce_SW2.r_CountZ0Z_0 ));
    Odrv4 I__1244 (
            .O(N__6423),
            .I(\Debounce_SW2.r_CountZ0Z_0 ));
    LocalMux I__1243 (
            .O(N__6420),
            .I(\Debounce_SW2.r_CountZ0Z_0 ));
    SRMux I__1242 (
            .O(N__6413),
            .I(N__6401));
    SRMux I__1241 (
            .O(N__6412),
            .I(N__6401));
    SRMux I__1240 (
            .O(N__6411),
            .I(N__6401));
    SRMux I__1239 (
            .O(N__6410),
            .I(N__6401));
    GlobalMux I__1238 (
            .O(N__6401),
            .I(N__6398));
    gio2CtrlBuf I__1237 (
            .O(N__6398),
            .I(\Debounce_SW2.N_38_g ));
    InMux I__1236 (
            .O(N__6395),
            .I(N__6387));
    InMux I__1235 (
            .O(N__6394),
            .I(N__6387));
    InMux I__1234 (
            .O(N__6393),
            .I(N__6384));
    InMux I__1233 (
            .O(N__6392),
            .I(N__6381));
    LocalMux I__1232 (
            .O(N__6387),
            .I(\Debounce_SW3.r_CountZ0Z_0 ));
    LocalMux I__1231 (
            .O(N__6384),
            .I(\Debounce_SW3.r_CountZ0Z_0 ));
    LocalMux I__1230 (
            .O(N__6381),
            .I(\Debounce_SW3.r_CountZ0Z_0 ));
    CascadeMux I__1229 (
            .O(N__6374),
            .I(N__6370));
    InMux I__1228 (
            .O(N__6373),
            .I(N__6366));
    InMux I__1227 (
            .O(N__6370),
            .I(N__6363));
    InMux I__1226 (
            .O(N__6369),
            .I(N__6360));
    LocalMux I__1225 (
            .O(N__6366),
            .I(\Debounce_SW3.r_CountZ0Z_1 ));
    LocalMux I__1224 (
            .O(N__6363),
            .I(\Debounce_SW3.r_CountZ0Z_1 ));
    LocalMux I__1223 (
            .O(N__6360),
            .I(\Debounce_SW3.r_CountZ0Z_1 ));
    InMux I__1222 (
            .O(N__6353),
            .I(N__6349));
    InMux I__1221 (
            .O(N__6352),
            .I(N__6346));
    LocalMux I__1220 (
            .O(N__6349),
            .I(\Debounce_SW3.r_CountZ0Z_2 ));
    LocalMux I__1219 (
            .O(N__6346),
            .I(\Debounce_SW3.r_CountZ0Z_2 ));
    InMux I__1218 (
            .O(N__6341),
            .I(\Debounce_SW3.un2_r_count_cry_1 ));
    CascadeMux I__1217 (
            .O(N__6338),
            .I(N__6334));
    InMux I__1216 (
            .O(N__6337),
            .I(N__6331));
    InMux I__1215 (
            .O(N__6334),
            .I(N__6328));
    LocalMux I__1214 (
            .O(N__6331),
            .I(\Debounce_SW3.r_CountZ0Z_3 ));
    LocalMux I__1213 (
            .O(N__6328),
            .I(\Debounce_SW3.r_CountZ0Z_3 ));
    InMux I__1212 (
            .O(N__6323),
            .I(\Debounce_SW3.un2_r_count_cry_2 ));
    InMux I__1211 (
            .O(N__6320),
            .I(N__6317));
    LocalMux I__1210 (
            .O(N__6317),
            .I(N__6313));
    InMux I__1209 (
            .O(N__6316),
            .I(N__6310));
    Odrv4 I__1208 (
            .O(N__6313),
            .I(\Game_Inst.w_LFSR_Data_5 ));
    LocalMux I__1207 (
            .O(N__6310),
            .I(\Game_Inst.w_LFSR_Data_5 ));
    InMux I__1206 (
            .O(N__6305),
            .I(N__6302));
    LocalMux I__1205 (
            .O(N__6302),
            .I(N__6298));
    InMux I__1204 (
            .O(N__6301),
            .I(N__6295));
    Odrv4 I__1203 (
            .O(N__6298),
            .I(\Game_Inst.w_LFSR_Data_3 ));
    LocalMux I__1202 (
            .O(N__6295),
            .I(\Game_Inst.w_LFSR_Data_3 ));
    InMux I__1201 (
            .O(N__6290),
            .I(N__6287));
    LocalMux I__1200 (
            .O(N__6287),
            .I(N__6283));
    InMux I__1199 (
            .O(N__6286),
            .I(N__6280));
    Odrv4 I__1198 (
            .O(N__6283),
            .I(\Game_Inst.w_LFSR_Data_4 ));
    LocalMux I__1197 (
            .O(N__6280),
            .I(\Game_Inst.w_LFSR_Data_4 ));
    CascadeMux I__1196 (
            .O(N__6275),
            .I(\Debounce_SW2.N_183_cascade_ ));
    IoInMux I__1195 (
            .O(N__6272),
            .I(N__6269));
    LocalMux I__1194 (
            .O(N__6269),
            .I(N__6266));
    Span4Mux_s3_v I__1193 (
            .O(N__6266),
            .I(N__6263));
    Odrv4 I__1192 (
            .O(N__6263),
            .I(\Debounce_SW2.N_38 ));
    InMux I__1191 (
            .O(N__6260),
            .I(N__6256));
    InMux I__1190 (
            .O(N__6259),
            .I(N__6253));
    LocalMux I__1189 (
            .O(N__6256),
            .I(\Debounce_SW2.r_CountZ0Z_10 ));
    LocalMux I__1188 (
            .O(N__6253),
            .I(\Debounce_SW2.r_CountZ0Z_10 ));
    InMux I__1187 (
            .O(N__6248),
            .I(N__6244));
    InMux I__1186 (
            .O(N__6247),
            .I(N__6241));
    LocalMux I__1185 (
            .O(N__6244),
            .I(\Debounce_SW2.r_CountZ0Z_9 ));
    LocalMux I__1184 (
            .O(N__6241),
            .I(\Debounce_SW2.r_CountZ0Z_9 ));
    CascadeMux I__1183 (
            .O(N__6236),
            .I(N__6232));
    InMux I__1182 (
            .O(N__6235),
            .I(N__6229));
    InMux I__1181 (
            .O(N__6232),
            .I(N__6226));
    LocalMux I__1180 (
            .O(N__6229),
            .I(\Debounce_SW2.r_CountZ0Z_11 ));
    LocalMux I__1179 (
            .O(N__6226),
            .I(\Debounce_SW2.r_CountZ0Z_11 ));
    InMux I__1178 (
            .O(N__6221),
            .I(N__6217));
    InMux I__1177 (
            .O(N__6220),
            .I(N__6214));
    LocalMux I__1176 (
            .O(N__6217),
            .I(\Debounce_SW2.r_CountZ0Z_8 ));
    LocalMux I__1175 (
            .O(N__6214),
            .I(\Debounce_SW2.r_CountZ0Z_8 ));
    CascadeMux I__1174 (
            .O(N__6209),
            .I(N__6204));
    InMux I__1173 (
            .O(N__6208),
            .I(N__6201));
    InMux I__1172 (
            .O(N__6207),
            .I(N__6198));
    InMux I__1171 (
            .O(N__6204),
            .I(N__6195));
    LocalMux I__1170 (
            .O(N__6201),
            .I(\Debounce_SW2.r_CountZ0Z_13 ));
    LocalMux I__1169 (
            .O(N__6198),
            .I(\Debounce_SW2.r_CountZ0Z_13 ));
    LocalMux I__1168 (
            .O(N__6195),
            .I(\Debounce_SW2.r_CountZ0Z_13 ));
    InMux I__1167 (
            .O(N__6188),
            .I(N__6183));
    InMux I__1166 (
            .O(N__6187),
            .I(N__6178));
    InMux I__1165 (
            .O(N__6186),
            .I(N__6178));
    LocalMux I__1164 (
            .O(N__6183),
            .I(\Debounce_SW2.r_CountZ0Z_12 ));
    LocalMux I__1163 (
            .O(N__6178),
            .I(\Debounce_SW2.r_CountZ0Z_12 ));
    CascadeMux I__1162 (
            .O(N__6173),
            .I(\Debounce_SW2.un9_r_count_0_a2_2_cascade_ ));
    InMux I__1161 (
            .O(N__6170),
            .I(N__6164));
    InMux I__1160 (
            .O(N__6169),
            .I(N__6164));
    LocalMux I__1159 (
            .O(N__6164),
            .I(\Debounce_SW2.N_160 ));
    InMux I__1158 (
            .O(N__6161),
            .I(N__6157));
    InMux I__1157 (
            .O(N__6160),
            .I(N__6154));
    LocalMux I__1156 (
            .O(N__6157),
            .I(\Debounce_SW2.r_CountZ0Z_6 ));
    LocalMux I__1155 (
            .O(N__6154),
            .I(\Debounce_SW2.r_CountZ0Z_6 ));
    InMux I__1154 (
            .O(N__6149),
            .I(N__6145));
    InMux I__1153 (
            .O(N__6148),
            .I(N__6142));
    LocalMux I__1152 (
            .O(N__6145),
            .I(\Debounce_SW2.r_CountZ0Z_5 ));
    LocalMux I__1151 (
            .O(N__6142),
            .I(\Debounce_SW2.r_CountZ0Z_5 ));
    InMux I__1150 (
            .O(N__6137),
            .I(N__6133));
    InMux I__1149 (
            .O(N__6136),
            .I(N__6130));
    LocalMux I__1148 (
            .O(N__6133),
            .I(\Debounce_SW2.r_CountZ0Z_4 ));
    LocalMux I__1147 (
            .O(N__6130),
            .I(\Debounce_SW2.r_CountZ0Z_4 ));
    CascadeMux I__1146 (
            .O(N__6125),
            .I(N__6122));
    InMux I__1145 (
            .O(N__6122),
            .I(N__6119));
    LocalMux I__1144 (
            .O(N__6119),
            .I(\Debounce_SW2.N_147 ));
    InMux I__1143 (
            .O(N__6116),
            .I(N__6113));
    LocalMux I__1142 (
            .O(N__6113),
            .I(\Game_Inst.r_Pattern_4Z0Z_1 ));
    InMux I__1141 (
            .O(N__6110),
            .I(N__6107));
    LocalMux I__1140 (
            .O(N__6107),
            .I(\Game_Inst.r_Pattern_4Z0Z_0 ));
    InMux I__1139 (
            .O(N__6104),
            .I(N__6101));
    LocalMux I__1138 (
            .O(N__6101),
            .I(N__6098));
    Span4Mux_h I__1137 (
            .O(N__6098),
            .I(N__6094));
    InMux I__1136 (
            .O(N__6097),
            .I(N__6091));
    Odrv4 I__1135 (
            .O(N__6094),
            .I(\Game_Inst.w_LFSR_Data_15 ));
    LocalMux I__1134 (
            .O(N__6091),
            .I(\Game_Inst.w_LFSR_Data_15 ));
    InMux I__1133 (
            .O(N__6086),
            .I(N__6083));
    LocalMux I__1132 (
            .O(N__6083),
            .I(\Game_Inst.r_Pattern_7Z0Z_1 ));
    InMux I__1131 (
            .O(N__6080),
            .I(N__6077));
    LocalMux I__1130 (
            .O(N__6077),
            .I(\Game_Inst.r_Pattern_5Z0Z_1 ));
    CEMux I__1129 (
            .O(N__6074),
            .I(N__6071));
    LocalMux I__1128 (
            .O(N__6071),
            .I(N__6068));
    Span4Mux_v I__1127 (
            .O(N__6068),
            .I(N__6063));
    CEMux I__1126 (
            .O(N__6067),
            .I(N__6060));
    CEMux I__1125 (
            .O(N__6066),
            .I(N__6057));
    Span4Mux_s3_h I__1124 (
            .O(N__6063),
            .I(N__6052));
    LocalMux I__1123 (
            .O(N__6060),
            .I(N__6052));
    LocalMux I__1122 (
            .O(N__6057),
            .I(N__6049));
    Odrv4 I__1121 (
            .O(N__6052),
            .I(\Game_Inst.r_SM_Main_d_6 ));
    Odrv4 I__1120 (
            .O(N__6049),
            .I(\Game_Inst.r_SM_Main_d_6 ));
    InMux I__1119 (
            .O(N__6044),
            .I(N__6037));
    InMux I__1118 (
            .O(N__6043),
            .I(N__6037));
    InMux I__1117 (
            .O(N__6042),
            .I(N__6034));
    LocalMux I__1116 (
            .O(N__6037),
            .I(N_143));
    LocalMux I__1115 (
            .O(N__6034),
            .I(N_143));
    InMux I__1114 (
            .O(N__6029),
            .I(N__6026));
    LocalMux I__1113 (
            .O(N__6026),
            .I(N__6022));
    InMux I__1112 (
            .O(N__6025),
            .I(N__6019));
    Odrv4 I__1111 (
            .O(N__6022),
            .I(\Game_Inst.w_LFSR_Data_7 ));
    LocalMux I__1110 (
            .O(N__6019),
            .I(\Game_Inst.w_LFSR_Data_7 ));
    InMux I__1109 (
            .O(N__6014),
            .I(N__6010));
    InMux I__1108 (
            .O(N__6013),
            .I(N__6007));
    LocalMux I__1107 (
            .O(N__6010),
            .I(N__6004));
    LocalMux I__1106 (
            .O(N__6007),
            .I(\Game_Inst.w_LFSR_Data_2 ));
    Odrv4 I__1105 (
            .O(N__6004),
            .I(\Game_Inst.w_LFSR_Data_2 ));
    InMux I__1104 (
            .O(N__5999),
            .I(N__5995));
    InMux I__1103 (
            .O(N__5998),
            .I(N__5992));
    LocalMux I__1102 (
            .O(N__5995),
            .I(\Game_Inst.w_LFSR_Data_6 ));
    LocalMux I__1101 (
            .O(N__5992),
            .I(\Game_Inst.w_LFSR_Data_6 ));
    CascadeMux I__1100 (
            .O(N__5987),
            .I(\Game_Inst.N_208_cascade_ ));
    InMux I__1099 (
            .O(N__5984),
            .I(N__5981));
    LocalMux I__1098 (
            .O(N__5981),
            .I(\Game_Inst.N_264 ));
    InMux I__1097 (
            .O(N__5978),
            .I(N__5975));
    LocalMux I__1096 (
            .O(N__5975),
            .I(\Game_Inst.r_Pattern_5Z0Z_0 ));
    InMux I__1095 (
            .O(N__5972),
            .I(N__5969));
    LocalMux I__1094 (
            .O(N__5969),
            .I(\Game_Inst.r_Pattern_3Z0Z_1 ));
    InMux I__1093 (
            .O(N__5966),
            .I(N__5963));
    LocalMux I__1092 (
            .O(N__5963),
            .I(\Game_Inst.r_Pattern_2Z0Z_1 ));
    InMux I__1091 (
            .O(N__5960),
            .I(N__5956));
    InMux I__1090 (
            .O(N__5959),
            .I(N__5953));
    LocalMux I__1089 (
            .O(N__5956),
            .I(N__5950));
    LocalMux I__1088 (
            .O(N__5953),
            .I(N__5947));
    Span4Mux_h I__1087 (
            .O(N__5950),
            .I(N__5944));
    Span4Mux_v I__1086 (
            .O(N__5947),
            .I(N__5941));
    Odrv4 I__1085 (
            .O(N__5944),
            .I(\Game_Inst.w_LFSR_Data_1 ));
    Odrv4 I__1084 (
            .O(N__5941),
            .I(\Game_Inst.w_LFSR_Data_1 ));
    InMux I__1083 (
            .O(N__5936),
            .I(N__5933));
    LocalMux I__1082 (
            .O(N__5933),
            .I(N__5930));
    Odrv4 I__1081 (
            .O(N__5930),
            .I(\Game_Inst.r_Pattern_0Z0Z_1 ));
    InMux I__1080 (
            .O(N__5927),
            .I(N__5924));
    LocalMux I__1079 (
            .O(N__5924),
            .I(\Game_Inst.r_Pattern_1Z0Z_1 ));
    InMux I__1078 (
            .O(N__5921),
            .I(N__5918));
    LocalMux I__1077 (
            .O(N__5918),
            .I(\Game_Inst.r_Pattern_6Z0Z_1 ));
    InMux I__1076 (
            .O(N__5915),
            .I(N__5912));
    LocalMux I__1075 (
            .O(N__5912),
            .I(\Game_Inst.r_Pattern_2Z0Z_0 ));
    InMux I__1074 (
            .O(N__5909),
            .I(N__5906));
    LocalMux I__1073 (
            .O(N__5906),
            .I(\Game_Inst.r_Pattern_3Z0Z_0 ));
    CascadeMux I__1072 (
            .O(N__5903),
            .I(N__5900));
    InMux I__1071 (
            .O(N__5900),
            .I(N__5896));
    InMux I__1070 (
            .O(N__5899),
            .I(N__5892));
    LocalMux I__1069 (
            .O(N__5896),
            .I(N__5889));
    InMux I__1068 (
            .O(N__5895),
            .I(N__5886));
    LocalMux I__1067 (
            .O(N__5892),
            .I(\Debounce_SW1.r_CountZ0Z_1 ));
    Odrv12 I__1066 (
            .O(N__5889),
            .I(\Debounce_SW1.r_CountZ0Z_1 ));
    LocalMux I__1065 (
            .O(N__5886),
            .I(\Debounce_SW1.r_CountZ0Z_1 ));
    InMux I__1064 (
            .O(N__5879),
            .I(N__5874));
    InMux I__1063 (
            .O(N__5878),
            .I(N__5868));
    InMux I__1062 (
            .O(N__5877),
            .I(N__5868));
    LocalMux I__1061 (
            .O(N__5874),
            .I(N__5865));
    InMux I__1060 (
            .O(N__5873),
            .I(N__5862));
    LocalMux I__1059 (
            .O(N__5868),
            .I(\Debounce_SW1.r_CountZ0Z_0 ));
    Odrv12 I__1058 (
            .O(N__5865),
            .I(\Debounce_SW1.r_CountZ0Z_0 ));
    LocalMux I__1057 (
            .O(N__5862),
            .I(\Debounce_SW1.r_CountZ0Z_0 ));
    SRMux I__1056 (
            .O(N__5855),
            .I(N__5843));
    SRMux I__1055 (
            .O(N__5854),
            .I(N__5843));
    SRMux I__1054 (
            .O(N__5853),
            .I(N__5843));
    SRMux I__1053 (
            .O(N__5852),
            .I(N__5843));
    GlobalMux I__1052 (
            .O(N__5843),
            .I(N__5840));
    gio2CtrlBuf I__1051 (
            .O(N__5840),
            .I(\Debounce_SW1.N_36_g ));
    InMux I__1050 (
            .O(N__5837),
            .I(N__5833));
    InMux I__1049 (
            .O(N__5836),
            .I(N__5830));
    LocalMux I__1048 (
            .O(N__5833),
            .I(N__5827));
    LocalMux I__1047 (
            .O(N__5830),
            .I(N__5824));
    Span4Mux_v I__1046 (
            .O(N__5827),
            .I(N__5821));
    Span4Mux_v I__1045 (
            .O(N__5824),
            .I(N__5818));
    Odrv4 I__1044 (
            .O(N__5821),
            .I(\Debounce_SW1.N_146 ));
    Odrv4 I__1043 (
            .O(N__5818),
            .I(\Debounce_SW1.N_146 ));
    InMux I__1042 (
            .O(N__5813),
            .I(N__5808));
    InMux I__1041 (
            .O(N__5812),
            .I(N__5805));
    InMux I__1040 (
            .O(N__5811),
            .I(N__5802));
    LocalMux I__1039 (
            .O(N__5808),
            .I(N__5799));
    LocalMux I__1038 (
            .O(N__5805),
            .I(N__5796));
    LocalMux I__1037 (
            .O(N__5802),
            .I(\Debounce_SW1.r_CountZ0Z_12 ));
    Odrv12 I__1036 (
            .O(N__5799),
            .I(\Debounce_SW1.r_CountZ0Z_12 ));
    Odrv4 I__1035 (
            .O(N__5796),
            .I(\Debounce_SW1.r_CountZ0Z_12 ));
    CascadeMux I__1034 (
            .O(N__5789),
            .I(N__5786));
    InMux I__1033 (
            .O(N__5786),
            .I(N__5783));
    LocalMux I__1032 (
            .O(N__5783),
            .I(N__5778));
    InMux I__1031 (
            .O(N__5782),
            .I(N__5775));
    InMux I__1030 (
            .O(N__5781),
            .I(N__5772));
    Span4Mux_h I__1029 (
            .O(N__5778),
            .I(N__5767));
    LocalMux I__1028 (
            .O(N__5775),
            .I(N__5767));
    LocalMux I__1027 (
            .O(N__5772),
            .I(\Debounce_SW1.r_CountZ0Z_13 ));
    Odrv4 I__1026 (
            .O(N__5767),
            .I(\Debounce_SW1.r_CountZ0Z_13 ));
    InMux I__1025 (
            .O(N__5762),
            .I(N__5758));
    InMux I__1024 (
            .O(N__5761),
            .I(N__5755));
    LocalMux I__1023 (
            .O(N__5758),
            .I(N__5749));
    LocalMux I__1022 (
            .O(N__5755),
            .I(N__5749));
    InMux I__1021 (
            .O(N__5754),
            .I(N__5746));
    Span4Mux_h I__1020 (
            .O(N__5749),
            .I(N__5743));
    LocalMux I__1019 (
            .O(N__5746),
            .I(\Debounce_SW1.r_CountZ0Z_7 ));
    Odrv4 I__1018 (
            .O(N__5743),
            .I(\Debounce_SW1.r_CountZ0Z_7 ));
    InMux I__1017 (
            .O(N__5738),
            .I(N__5735));
    LocalMux I__1016 (
            .O(N__5735),
            .I(\Debounce_SW1.un9_r_count_10 ));
    InMux I__1015 (
            .O(N__5732),
            .I(N__5729));
    LocalMux I__1014 (
            .O(N__5729),
            .I(N__5725));
    InMux I__1013 (
            .O(N__5728),
            .I(N__5722));
    Span4Mux_h I__1012 (
            .O(N__5725),
            .I(N__5717));
    LocalMux I__1011 (
            .O(N__5722),
            .I(N__5717));
    Odrv4 I__1010 (
            .O(N__5717),
            .I(\Debounce_SW1.r_count15_i_a2_0 ));
    CascadeMux I__1009 (
            .O(N__5714),
            .I(\Debounce_SW1.un9_r_count_0_a2_2_cascade_ ));
    InMux I__1008 (
            .O(N__5711),
            .I(N__5707));
    InMux I__1007 (
            .O(N__5710),
            .I(N__5704));
    LocalMux I__1006 (
            .O(N__5707),
            .I(N__5699));
    LocalMux I__1005 (
            .O(N__5704),
            .I(N__5699));
    Odrv12 I__1004 (
            .O(N__5699),
            .I(\Debounce_SW1.N_161 ));
    InMux I__1003 (
            .O(N__5696),
            .I(N__5693));
    LocalMux I__1002 (
            .O(N__5693),
            .I(\Game_Inst.r_SwitchZ0Z_4 ));
    InMux I__1001 (
            .O(N__5690),
            .I(N__5687));
    LocalMux I__1000 (
            .O(N__5687),
            .I(\Game_Inst.r_SwitchZ0Z_2 ));
    InMux I__999 (
            .O(N__5684),
            .I(N__5675));
    InMux I__998 (
            .O(N__5683),
            .I(N__5675));
    InMux I__997 (
            .O(N__5682),
            .I(N__5675));
    LocalMux I__996 (
            .O(N__5675),
            .I(\Game_Inst.r_Switch_1_RNIA12HZ0 ));
    InMux I__995 (
            .O(N__5672),
            .I(N__5669));
    LocalMux I__994 (
            .O(N__5669),
            .I(\Game_Inst.r_SwitchZ0Z_1 ));
    CascadeMux I__993 (
            .O(N__5666),
            .I(N__5662));
    CascadeMux I__992 (
            .O(N__5665),
            .I(N__5658));
    InMux I__991 (
            .O(N__5662),
            .I(N__5652));
    InMux I__990 (
            .O(N__5661),
            .I(N__5652));
    InMux I__989 (
            .O(N__5658),
            .I(N__5649));
    InMux I__988 (
            .O(N__5657),
            .I(N__5644));
    LocalMux I__987 (
            .O(N__5652),
            .I(N__5640));
    LocalMux I__986 (
            .O(N__5649),
            .I(N__5637));
    CascadeMux I__985 (
            .O(N__5648),
            .I(N__5634));
    InMux I__984 (
            .O(N__5647),
            .I(N__5631));
    LocalMux I__983 (
            .O(N__5644),
            .I(N__5628));
    InMux I__982 (
            .O(N__5643),
            .I(N__5625));
    Span4Mux_v I__981 (
            .O(N__5640),
            .I(N__5620));
    Span4Mux_v I__980 (
            .O(N__5637),
            .I(N__5620));
    InMux I__979 (
            .O(N__5634),
            .I(N__5617));
    LocalMux I__978 (
            .O(N__5631),
            .I(N__5612));
    Span4Mux_h I__977 (
            .O(N__5628),
            .I(N__5612));
    LocalMux I__976 (
            .O(N__5625),
            .I(\Game_Inst.w_Toggle ));
    Odrv4 I__975 (
            .O(N__5620),
            .I(\Game_Inst.w_Toggle ));
    LocalMux I__974 (
            .O(N__5617),
            .I(\Game_Inst.w_Toggle ));
    Odrv4 I__973 (
            .O(N__5612),
            .I(\Game_Inst.w_Toggle ));
    InMux I__972 (
            .O(N__5603),
            .I(N__5594));
    InMux I__971 (
            .O(N__5602),
            .I(N__5594));
    InMux I__970 (
            .O(N__5601),
            .I(N__5594));
    LocalMux I__969 (
            .O(N__5594),
            .I(N__5589));
    InMux I__968 (
            .O(N__5593),
            .I(N__5586));
    InMux I__967 (
            .O(N__5592),
            .I(N__5583));
    Odrv4 I__966 (
            .O(N__5589),
            .I(\Game_Inst.r_ToggleZ0 ));
    LocalMux I__965 (
            .O(N__5586),
            .I(\Game_Inst.r_ToggleZ0 ));
    LocalMux I__964 (
            .O(N__5583),
            .I(\Game_Inst.r_ToggleZ0 ));
    InMux I__963 (
            .O(N__5576),
            .I(N__5573));
    LocalMux I__962 (
            .O(N__5573),
            .I(\Debounce_SW3.N_159 ));
    CascadeMux I__961 (
            .O(N__5570),
            .I(\Debounce_SW3.N_159_cascade_ ));
    InMux I__960 (
            .O(N__5567),
            .I(N__5564));
    LocalMux I__959 (
            .O(N__5564),
            .I(\Debounce_SW3.N_287 ));
    InMux I__958 (
            .O(N__5561),
            .I(N__5558));
    LocalMux I__957 (
            .O(N__5558),
            .I(\Debounce_SW3.un9_r_count_0_a2_2 ));
    InMux I__956 (
            .O(N__5555),
            .I(N__5549));
    InMux I__955 (
            .O(N__5554),
            .I(N__5549));
    LocalMux I__954 (
            .O(N__5549),
            .I(\Debounce_SW3.N_148 ));
    CascadeMux I__953 (
            .O(N__5546),
            .I(\Debounce_SW3.r_count15_i_a2_0_cascade_ ));
    InMux I__952 (
            .O(N__5543),
            .I(N__5537));
    InMux I__951 (
            .O(N__5542),
            .I(N__5537));
    LocalMux I__950 (
            .O(N__5537),
            .I(\Debounce_SW3.un9_r_count_10 ));
    InMux I__949 (
            .O(N__5534),
            .I(N__5530));
    InMux I__948 (
            .O(N__5533),
            .I(N__5527));
    LocalMux I__947 (
            .O(N__5530),
            .I(\Debounce_SW4.r_CountZ0Z_15 ));
    LocalMux I__946 (
            .O(N__5527),
            .I(\Debounce_SW4.r_CountZ0Z_15 ));
    InMux I__945 (
            .O(N__5522),
            .I(N__5518));
    InMux I__944 (
            .O(N__5521),
            .I(N__5515));
    LocalMux I__943 (
            .O(N__5518),
            .I(N__5512));
    LocalMux I__942 (
            .O(N__5515),
            .I(\Debounce_SW4.r_CountZ0Z_16 ));
    Odrv4 I__941 (
            .O(N__5512),
            .I(\Debounce_SW4.r_CountZ0Z_16 ));
    CascadeMux I__940 (
            .O(N__5507),
            .I(N__5504));
    InMux I__939 (
            .O(N__5504),
            .I(N__5501));
    LocalMux I__938 (
            .O(N__5501),
            .I(N__5497));
    InMux I__937 (
            .O(N__5500),
            .I(N__5494));
    Span4Mux_h I__936 (
            .O(N__5497),
            .I(N__5491));
    LocalMux I__935 (
            .O(N__5494),
            .I(\Debounce_SW4.r_CountZ0Z_14 ));
    Odrv4 I__934 (
            .O(N__5491),
            .I(\Debounce_SW4.r_CountZ0Z_14 ));
    InMux I__933 (
            .O(N__5486),
            .I(N__5482));
    InMux I__932 (
            .O(N__5485),
            .I(N__5479));
    LocalMux I__931 (
            .O(N__5482),
            .I(\Debounce_SW4.r_CountZ0Z_17 ));
    LocalMux I__930 (
            .O(N__5479),
            .I(\Debounce_SW4.r_CountZ0Z_17 ));
    InMux I__929 (
            .O(N__5474),
            .I(N__5470));
    InMux I__928 (
            .O(N__5473),
            .I(N__5467));
    LocalMux I__927 (
            .O(N__5470),
            .I(N__5464));
    LocalMux I__926 (
            .O(N__5467),
            .I(N__5459));
    Span4Mux_s2_v I__925 (
            .O(N__5464),
            .I(N__5459));
    Odrv4 I__924 (
            .O(N__5459),
            .I(\Debounce_SW4.r_count15_i_a2_0 ));
    InMux I__923 (
            .O(N__5456),
            .I(\Debounce_SW2.un2_r_count_cry_11 ));
    InMux I__922 (
            .O(N__5453),
            .I(\Debounce_SW2.un2_r_count_cry_12 ));
    InMux I__921 (
            .O(N__5450),
            .I(\Debounce_SW2.un2_r_count_cry_13 ));
    InMux I__920 (
            .O(N__5447),
            .I(\Debounce_SW2.un2_r_count_cry_14 ));
    InMux I__919 (
            .O(N__5444),
            .I(\Debounce_SW2.un2_r_count_cry_15 ));
    InMux I__918 (
            .O(N__5441),
            .I(bfn_7_15_0_));
    InMux I__917 (
            .O(N__5438),
            .I(N__5435));
    LocalMux I__916 (
            .O(N__5435),
            .I(N__5431));
    InMux I__915 (
            .O(N__5434),
            .I(N__5428));
    Span4Mux_s3_v I__914 (
            .O(N__5431),
            .I(N__5425));
    LocalMux I__913 (
            .O(N__5428),
            .I(N__5422));
    Span4Mux_h I__912 (
            .O(N__5425),
            .I(N__5419));
    Span4Mux_s3_v I__911 (
            .O(N__5422),
            .I(N__5416));
    Odrv4 I__910 (
            .O(N__5419),
            .I(i_Switch_4_c));
    Odrv4 I__909 (
            .O(N__5416),
            .I(i_Switch_4_c));
    CEMux I__908 (
            .O(N__5411),
            .I(N__5408));
    LocalMux I__907 (
            .O(N__5408),
            .I(N__5405));
    Odrv4 I__906 (
            .O(N__5405),
            .I(\Debounce_SW4.r_State_e_0_RNO_2 ));
    InMux I__905 (
            .O(N__5402),
            .I(\Debounce_SW2.un2_r_count_cry_2 ));
    InMux I__904 (
            .O(N__5399),
            .I(\Debounce_SW2.un2_r_count_cry_3 ));
    InMux I__903 (
            .O(N__5396),
            .I(\Debounce_SW2.un2_r_count_cry_4 ));
    InMux I__902 (
            .O(N__5393),
            .I(\Debounce_SW2.un2_r_count_cry_5 ));
    InMux I__901 (
            .O(N__5390),
            .I(\Debounce_SW2.un2_r_count_cry_6 ));
    InMux I__900 (
            .O(N__5387),
            .I(\Debounce_SW2.un2_r_count_cry_7 ));
    InMux I__899 (
            .O(N__5384),
            .I(bfn_7_14_0_));
    InMux I__898 (
            .O(N__5381),
            .I(\Debounce_SW2.un2_r_count_cry_9 ));
    InMux I__897 (
            .O(N__5378),
            .I(\Debounce_SW2.un2_r_count_cry_10 ));
    InMux I__896 (
            .O(N__5375),
            .I(N__5372));
    LocalMux I__895 (
            .O(N__5372),
            .I(N__5368));
    InMux I__894 (
            .O(N__5371),
            .I(N__5365));
    Span4Mux_h I__893 (
            .O(N__5368),
            .I(N__5358));
    LocalMux I__892 (
            .O(N__5365),
            .I(N__5358));
    InMux I__891 (
            .O(N__5364),
            .I(N__5353));
    InMux I__890 (
            .O(N__5363),
            .I(N__5353));
    Odrv4 I__889 (
            .O(N__5358),
            .I(\Game_Inst.r_Button_DVZ0 ));
    LocalMux I__888 (
            .O(N__5353),
            .I(\Game_Inst.r_Button_DVZ0 ));
    CascadeMux I__887 (
            .O(N__5348),
            .I(\Game_Inst.r_SM_Main_d_6_cascade_ ));
    CascadeMux I__886 (
            .O(N__5345),
            .I(N__5341));
    InMux I__885 (
            .O(N__5344),
            .I(N__5323));
    InMux I__884 (
            .O(N__5341),
            .I(N__5323));
    InMux I__883 (
            .O(N__5340),
            .I(N__5323));
    InMux I__882 (
            .O(N__5339),
            .I(N__5320));
    InMux I__881 (
            .O(N__5338),
            .I(N__5317));
    InMux I__880 (
            .O(N__5337),
            .I(N__5314));
    InMux I__879 (
            .O(N__5336),
            .I(N__5305));
    InMux I__878 (
            .O(N__5335),
            .I(N__5305));
    InMux I__877 (
            .O(N__5334),
            .I(N__5305));
    InMux I__876 (
            .O(N__5333),
            .I(N__5305));
    InMux I__875 (
            .O(N__5332),
            .I(N__5300));
    InMux I__874 (
            .O(N__5331),
            .I(N__5300));
    InMux I__873 (
            .O(N__5330),
            .I(N__5297));
    LocalMux I__872 (
            .O(N__5323),
            .I(\Game_Inst.r_IndexZ1Z_0 ));
    LocalMux I__871 (
            .O(N__5320),
            .I(\Game_Inst.r_IndexZ1Z_0 ));
    LocalMux I__870 (
            .O(N__5317),
            .I(\Game_Inst.r_IndexZ1Z_0 ));
    LocalMux I__869 (
            .O(N__5314),
            .I(\Game_Inst.r_IndexZ1Z_0 ));
    LocalMux I__868 (
            .O(N__5305),
            .I(\Game_Inst.r_IndexZ1Z_0 ));
    LocalMux I__867 (
            .O(N__5300),
            .I(\Game_Inst.r_IndexZ1Z_0 ));
    LocalMux I__866 (
            .O(N__5297),
            .I(\Game_Inst.r_IndexZ1Z_0 ));
    InMux I__865 (
            .O(N__5282),
            .I(N__5279));
    LocalMux I__864 (
            .O(N__5279),
            .I(N__5276));
    Odrv4 I__863 (
            .O(N__5276),
            .I(\Game_Inst.r_Pattern_4_RNILI2AZ0Z_0 ));
    InMux I__862 (
            .O(N__5273),
            .I(N__5270));
    LocalMux I__861 (
            .O(N__5270),
            .I(\Game_Inst.N_259 ));
    CascadeMux I__860 (
            .O(N__5267),
            .I(\Game_Inst.r_SM_Main_ns_i_0_1_2_cascade_ ));
    InMux I__859 (
            .O(N__5264),
            .I(N__5260));
    InMux I__858 (
            .O(N__5263),
            .I(N__5257));
    LocalMux I__857 (
            .O(N__5260),
            .I(\Game_Inst.N_260_1 ));
    LocalMux I__856 (
            .O(N__5257),
            .I(\Game_Inst.N_260_1 ));
    InMux I__855 (
            .O(N__5252),
            .I(\Debounce_SW2.un2_r_count_cry_1 ));
    InMux I__854 (
            .O(N__5249),
            .I(N__5241));
    InMux I__853 (
            .O(N__5248),
            .I(N__5238));
    InMux I__852 (
            .O(N__5247),
            .I(N__5231));
    InMux I__851 (
            .O(N__5246),
            .I(N__5231));
    InMux I__850 (
            .O(N__5245),
            .I(N__5231));
    InMux I__849 (
            .O(N__5244),
            .I(N__5228));
    LocalMux I__848 (
            .O(N__5241),
            .I(\Game_Inst.r_IndexZ0Z_1 ));
    LocalMux I__847 (
            .O(N__5238),
            .I(\Game_Inst.r_IndexZ0Z_1 ));
    LocalMux I__846 (
            .O(N__5231),
            .I(\Game_Inst.r_IndexZ0Z_1 ));
    LocalMux I__845 (
            .O(N__5228),
            .I(\Game_Inst.r_IndexZ0Z_1 ));
    CascadeMux I__844 (
            .O(N__5219),
            .I(\Game_Inst.r_Pattern_0_RNIFS911Z0Z_1_cascade_ ));
    InMux I__843 (
            .O(N__5216),
            .I(N__5208));
    InMux I__842 (
            .O(N__5215),
            .I(N__5201));
    InMux I__841 (
            .O(N__5214),
            .I(N__5201));
    InMux I__840 (
            .O(N__5213),
            .I(N__5201));
    InMux I__839 (
            .O(N__5212),
            .I(N__5196));
    InMux I__838 (
            .O(N__5211),
            .I(N__5196));
    LocalMux I__837 (
            .O(N__5208),
            .I(\Game_Inst.r_IndexZ0Z_2 ));
    LocalMux I__836 (
            .O(N__5201),
            .I(\Game_Inst.r_IndexZ0Z_2 ));
    LocalMux I__835 (
            .O(N__5196),
            .I(\Game_Inst.r_IndexZ0Z_2 ));
    CascadeMux I__834 (
            .O(N__5189),
            .I(\Game_Inst.un6_r_button_dv_7_i_m2_ns_1_1_cascade_ ));
    InMux I__833 (
            .O(N__5186),
            .I(N__5183));
    LocalMux I__832 (
            .O(N__5183),
            .I(\Game_Inst.r_Pattern_3_RNIH6MLZ0Z_0 ));
    InMux I__831 (
            .O(N__5180),
            .I(N__5177));
    LocalMux I__830 (
            .O(N__5177),
            .I(\Game_Inst.r_Pattern_3_RNIJ8MLZ0Z_1 ));
    CascadeMux I__829 (
            .O(N__5174),
            .I(N__5171));
    InMux I__828 (
            .O(N__5171),
            .I(N__5168));
    LocalMux I__827 (
            .O(N__5168),
            .I(N__5163));
    InMux I__826 (
            .O(N__5167),
            .I(N__5158));
    InMux I__825 (
            .O(N__5166),
            .I(N__5158));
    Odrv4 I__824 (
            .O(N__5163),
            .I(\Game_Inst.N_303 ));
    LocalMux I__823 (
            .O(N__5158),
            .I(\Game_Inst.N_303 ));
    InMux I__822 (
            .O(N__5153),
            .I(N__5150));
    LocalMux I__821 (
            .O(N__5150),
            .I(N__5147));
    Odrv4 I__820 (
            .O(N__5147),
            .I(\Game_Inst.r_SM_Main_ns_i_0_2_0 ));
    InMux I__819 (
            .O(N__5144),
            .I(N__5141));
    LocalMux I__818 (
            .O(N__5141),
            .I(\Game_Inst.r_Pattern_6_RNIR0FEZ0Z_1 ));
    InMux I__817 (
            .O(N__5138),
            .I(N__5135));
    LocalMux I__816 (
            .O(N__5135),
            .I(\Game_Inst.r_Pattern_4_RNINK2AZ0Z_1 ));
    InMux I__815 (
            .O(N__5132),
            .I(N__5129));
    LocalMux I__814 (
            .O(N__5129),
            .I(\Game_Inst.N_266 ));
    CascadeMux I__813 (
            .O(N__5126),
            .I(\Debounce_SW1.un9_r_count_10_cascade_ ));
    CascadeMux I__812 (
            .O(N__5123),
            .I(\Debounce_SW1.N_285_cascade_ ));
    CascadeMux I__811 (
            .O(N__5120),
            .I(\Debounce_SW1.N_184_cascade_ ));
    IoInMux I__810 (
            .O(N__5117),
            .I(N__5114));
    LocalMux I__809 (
            .O(N__5114),
            .I(N__5111));
    Odrv12 I__808 (
            .O(N__5111),
            .I(\Debounce_SW1.N_36 ));
    InMux I__807 (
            .O(N__5108),
            .I(N__5105));
    LocalMux I__806 (
            .O(N__5105),
            .I(\Game_Inst.r_Button_IDZ0Z_0 ));
    CascadeMux I__805 (
            .O(N__5102),
            .I(\Game_Inst.N_255_cascade_ ));
    InMux I__804 (
            .O(N__5099),
            .I(N__5090));
    InMux I__803 (
            .O(N__5098),
            .I(N__5090));
    InMux I__802 (
            .O(N__5097),
            .I(N__5090));
    LocalMux I__801 (
            .O(N__5090),
            .I(\Game_Inst.N_167 ));
    CascadeMux I__800 (
            .O(N__5087),
            .I(N__5083));
    InMux I__799 (
            .O(N__5086),
            .I(N__5078));
    InMux I__798 (
            .O(N__5083),
            .I(N__5078));
    LocalMux I__797 (
            .O(N__5078),
            .I(\Game_Inst.N_255 ));
    InMux I__796 (
            .O(N__5075),
            .I(N__5072));
    LocalMux I__795 (
            .O(N__5072),
            .I(\Game_Inst.r_Button_IDZ0Z_1 ));
    InMux I__794 (
            .O(N__5069),
            .I(N__5065));
    InMux I__793 (
            .O(N__5068),
            .I(N__5062));
    LocalMux I__792 (
            .O(N__5065),
            .I(N__5059));
    LocalMux I__791 (
            .O(N__5062),
            .I(\Debounce_SW4.r_CountZ0Z_10 ));
    Odrv12 I__790 (
            .O(N__5059),
            .I(\Debounce_SW4.r_CountZ0Z_10 ));
    InMux I__789 (
            .O(N__5054),
            .I(\Debounce_SW4.un2_r_count_cry_9 ));
    CascadeMux I__788 (
            .O(N__5051),
            .I(N__5048));
    InMux I__787 (
            .O(N__5048),
            .I(N__5044));
    InMux I__786 (
            .O(N__5047),
            .I(N__5041));
    LocalMux I__785 (
            .O(N__5044),
            .I(N__5038));
    LocalMux I__784 (
            .O(N__5041),
            .I(\Debounce_SW4.r_CountZ0Z_11 ));
    Odrv4 I__783 (
            .O(N__5038),
            .I(\Debounce_SW4.r_CountZ0Z_11 ));
    InMux I__782 (
            .O(N__5033),
            .I(\Debounce_SW4.un2_r_count_cry_10 ));
    InMux I__781 (
            .O(N__5030),
            .I(N__5025));
    InMux I__780 (
            .O(N__5029),
            .I(N__5022));
    InMux I__779 (
            .O(N__5028),
            .I(N__5019));
    LocalMux I__778 (
            .O(N__5025),
            .I(N__5014));
    LocalMux I__777 (
            .O(N__5022),
            .I(N__5014));
    LocalMux I__776 (
            .O(N__5019),
            .I(\Debounce_SW4.r_CountZ0Z_12 ));
    Odrv4 I__775 (
            .O(N__5014),
            .I(\Debounce_SW4.r_CountZ0Z_12 ));
    InMux I__774 (
            .O(N__5009),
            .I(\Debounce_SW4.un2_r_count_cry_11 ));
    CascadeMux I__773 (
            .O(N__5006),
            .I(N__5002));
    InMux I__772 (
            .O(N__5005),
            .I(N__4998));
    InMux I__771 (
            .O(N__5002),
            .I(N__4995));
    InMux I__770 (
            .O(N__5001),
            .I(N__4992));
    LocalMux I__769 (
            .O(N__4998),
            .I(N__4987));
    LocalMux I__768 (
            .O(N__4995),
            .I(N__4987));
    LocalMux I__767 (
            .O(N__4992),
            .I(\Debounce_SW4.r_CountZ0Z_13 ));
    Odrv4 I__766 (
            .O(N__4987),
            .I(\Debounce_SW4.r_CountZ0Z_13 ));
    InMux I__765 (
            .O(N__4982),
            .I(\Debounce_SW4.un2_r_count_cry_12 ));
    InMux I__764 (
            .O(N__4979),
            .I(\Debounce_SW4.un2_r_count_cry_13 ));
    InMux I__763 (
            .O(N__4976),
            .I(\Debounce_SW4.un2_r_count_cry_14 ));
    InMux I__762 (
            .O(N__4973),
            .I(\Debounce_SW4.un2_r_count_cry_15 ));
    InMux I__761 (
            .O(N__4970),
            .I(bfn_7_7_0_));
    SRMux I__760 (
            .O(N__4967),
            .I(N__4955));
    SRMux I__759 (
            .O(N__4966),
            .I(N__4955));
    SRMux I__758 (
            .O(N__4965),
            .I(N__4955));
    SRMux I__757 (
            .O(N__4964),
            .I(N__4955));
    GlobalMux I__756 (
            .O(N__4955),
            .I(N__4952));
    gio2CtrlBuf I__755 (
            .O(N__4952),
            .I(\Debounce_SW4.N_42_g ));
    InMux I__754 (
            .O(N__4949),
            .I(N__4946));
    LocalMux I__753 (
            .O(N__4946),
            .I(N__4942));
    InMux I__752 (
            .O(N__4945),
            .I(N__4939));
    Span4Mux_h I__751 (
            .O(N__4942),
            .I(N__4936));
    LocalMux I__750 (
            .O(N__4939),
            .I(\Debounce_SW1.r_CountZ0Z_2 ));
    Odrv4 I__749 (
            .O(N__4936),
            .I(\Debounce_SW1.r_CountZ0Z_2 ));
    CascadeMux I__748 (
            .O(N__4931),
            .I(N__4928));
    InMux I__747 (
            .O(N__4928),
            .I(N__4925));
    LocalMux I__746 (
            .O(N__4925),
            .I(N__4921));
    InMux I__745 (
            .O(N__4924),
            .I(N__4918));
    Span4Mux_h I__744 (
            .O(N__4921),
            .I(N__4915));
    LocalMux I__743 (
            .O(N__4918),
            .I(\Debounce_SW1.r_CountZ0Z_3 ));
    Odrv4 I__742 (
            .O(N__4915),
            .I(\Debounce_SW1.r_CountZ0Z_3 ));
    InMux I__741 (
            .O(N__4910),
            .I(N__4906));
    InMux I__740 (
            .O(N__4909),
            .I(N__4903));
    LocalMux I__739 (
            .O(N__4906),
            .I(\Debounce_SW4.r_CountZ0Z_2 ));
    LocalMux I__738 (
            .O(N__4903),
            .I(\Debounce_SW4.r_CountZ0Z_2 ));
    InMux I__737 (
            .O(N__4898),
            .I(\Debounce_SW4.un2_r_count_cry_1 ));
    CascadeMux I__736 (
            .O(N__4895),
            .I(N__4891));
    InMux I__735 (
            .O(N__4894),
            .I(N__4888));
    InMux I__734 (
            .O(N__4891),
            .I(N__4885));
    LocalMux I__733 (
            .O(N__4888),
            .I(\Debounce_SW4.r_CountZ0Z_3 ));
    LocalMux I__732 (
            .O(N__4885),
            .I(\Debounce_SW4.r_CountZ0Z_3 ));
    InMux I__731 (
            .O(N__4880),
            .I(\Debounce_SW4.un2_r_count_cry_2 ));
    InMux I__730 (
            .O(N__4877),
            .I(N__4873));
    InMux I__729 (
            .O(N__4876),
            .I(N__4870));
    LocalMux I__728 (
            .O(N__4873),
            .I(\Debounce_SW4.r_CountZ0Z_4 ));
    LocalMux I__727 (
            .O(N__4870),
            .I(\Debounce_SW4.r_CountZ0Z_4 ));
    InMux I__726 (
            .O(N__4865),
            .I(\Debounce_SW4.un2_r_count_cry_3 ));
    InMux I__725 (
            .O(N__4862),
            .I(N__4858));
    InMux I__724 (
            .O(N__4861),
            .I(N__4855));
    LocalMux I__723 (
            .O(N__4858),
            .I(\Debounce_SW4.r_CountZ0Z_5 ));
    LocalMux I__722 (
            .O(N__4855),
            .I(\Debounce_SW4.r_CountZ0Z_5 ));
    InMux I__721 (
            .O(N__4850),
            .I(\Debounce_SW4.un2_r_count_cry_4 ));
    InMux I__720 (
            .O(N__4847),
            .I(N__4843));
    InMux I__719 (
            .O(N__4846),
            .I(N__4840));
    LocalMux I__718 (
            .O(N__4843),
            .I(\Debounce_SW4.r_CountZ0Z_6 ));
    LocalMux I__717 (
            .O(N__4840),
            .I(\Debounce_SW4.r_CountZ0Z_6 ));
    InMux I__716 (
            .O(N__4835),
            .I(\Debounce_SW4.un2_r_count_cry_5 ));
    InMux I__715 (
            .O(N__4832),
            .I(N__4827));
    InMux I__714 (
            .O(N__4831),
            .I(N__4822));
    InMux I__713 (
            .O(N__4830),
            .I(N__4822));
    LocalMux I__712 (
            .O(N__4827),
            .I(\Debounce_SW4.r_CountZ0Z_7 ));
    LocalMux I__711 (
            .O(N__4822),
            .I(\Debounce_SW4.r_CountZ0Z_7 ));
    InMux I__710 (
            .O(N__4817),
            .I(\Debounce_SW4.un2_r_count_cry_6 ));
    InMux I__709 (
            .O(N__4814),
            .I(N__4810));
    InMux I__708 (
            .O(N__4813),
            .I(N__4807));
    LocalMux I__707 (
            .O(N__4810),
            .I(\Debounce_SW4.r_CountZ0Z_8 ));
    LocalMux I__706 (
            .O(N__4807),
            .I(\Debounce_SW4.r_CountZ0Z_8 ));
    InMux I__705 (
            .O(N__4802),
            .I(\Debounce_SW4.un2_r_count_cry_7 ));
    InMux I__704 (
            .O(N__4799),
            .I(N__4795));
    InMux I__703 (
            .O(N__4798),
            .I(N__4792));
    LocalMux I__702 (
            .O(N__4795),
            .I(N__4789));
    LocalMux I__701 (
            .O(N__4792),
            .I(\Debounce_SW4.r_CountZ0Z_9 ));
    Odrv4 I__700 (
            .O(N__4789),
            .I(\Debounce_SW4.r_CountZ0Z_9 ));
    InMux I__699 (
            .O(N__4784),
            .I(bfn_7_6_0_));
    CascadeMux I__698 (
            .O(N__4781),
            .I(\Debounce_SW4.N_181_cascade_ ));
    IoInMux I__697 (
            .O(N__4778),
            .I(N__4775));
    LocalMux I__696 (
            .O(N__4775),
            .I(N__4772));
    Odrv4 I__695 (
            .O(N__4772),
            .I(\Debounce_SW4.N_42 ));
    CascadeMux I__694 (
            .O(N__4769),
            .I(\Debounce_SW4.un9_r_count_10_cascade_ ));
    InMux I__693 (
            .O(N__4766),
            .I(N__4763));
    LocalMux I__692 (
            .O(N__4763),
            .I(\Debounce_SW4.N_288 ));
    InMux I__691 (
            .O(N__4760),
            .I(N__4757));
    LocalMux I__690 (
            .O(N__4757),
            .I(\Debounce_SW4.N_158 ));
    CascadeMux I__689 (
            .O(N__4754),
            .I(\Debounce_SW4.N_158_cascade_ ));
    InMux I__688 (
            .O(N__4751),
            .I(N__4745));
    InMux I__687 (
            .O(N__4750),
            .I(N__4745));
    LocalMux I__686 (
            .O(N__4745),
            .I(\Debounce_SW4.N_149 ));
    InMux I__685 (
            .O(N__4742),
            .I(N__4739));
    LocalMux I__684 (
            .O(N__4739),
            .I(\Debounce_SW4.un9_r_count_10 ));
    CascadeMux I__683 (
            .O(N__4736),
            .I(\Debounce_SW4.un9_r_count_0_a2_2_cascade_ ));
    InMux I__682 (
            .O(N__4733),
            .I(N__4725));
    InMux I__681 (
            .O(N__4732),
            .I(N__4725));
    InMux I__680 (
            .O(N__4731),
            .I(N__4722));
    InMux I__679 (
            .O(N__4730),
            .I(N__4719));
    LocalMux I__678 (
            .O(N__4725),
            .I(\Debounce_SW4.r_CountZ0Z_0 ));
    LocalMux I__677 (
            .O(N__4722),
            .I(\Debounce_SW4.r_CountZ0Z_0 ));
    LocalMux I__676 (
            .O(N__4719),
            .I(\Debounce_SW4.r_CountZ0Z_0 ));
    CascadeMux I__675 (
            .O(N__4712),
            .I(N__4708));
    InMux I__674 (
            .O(N__4711),
            .I(N__4704));
    InMux I__673 (
            .O(N__4708),
            .I(N__4701));
    InMux I__672 (
            .O(N__4707),
            .I(N__4698));
    LocalMux I__671 (
            .O(N__4704),
            .I(\Debounce_SW4.r_CountZ0Z_1 ));
    LocalMux I__670 (
            .O(N__4701),
            .I(\Debounce_SW4.r_CountZ0Z_1 ));
    LocalMux I__669 (
            .O(N__4698),
            .I(\Debounce_SW4.r_CountZ0Z_1 ));
    InMux I__668 (
            .O(N__4691),
            .I(N__4688));
    LocalMux I__667 (
            .O(N__4688),
            .I(\Game_Inst.r_Pattern_7Z0Z_0 ));
    InMux I__666 (
            .O(N__4685),
            .I(N__4682));
    LocalMux I__665 (
            .O(N__4682),
            .I(\Game_Inst.r_Pattern_6Z0Z_0 ));
    InMux I__664 (
            .O(N__4679),
            .I(N__4676));
    LocalMux I__663 (
            .O(N__4676),
            .I(N__4673));
    Odrv4 I__662 (
            .O(N__4673),
            .I(\Game_Inst.r_Pattern_6_RNIPUEEZ0Z_0 ));
    InMux I__661 (
            .O(N__4670),
            .I(N__4665));
    InMux I__660 (
            .O(N__4669),
            .I(N__4659));
    InMux I__659 (
            .O(N__4668),
            .I(N__4659));
    LocalMux I__658 (
            .O(N__4665),
            .I(N__4656));
    InMux I__657 (
            .O(N__4664),
            .I(N__4653));
    LocalMux I__656 (
            .O(N__4659),
            .I(\Game_Inst.N_132 ));
    Odrv4 I__655 (
            .O(N__4656),
            .I(\Game_Inst.N_132 ));
    LocalMux I__654 (
            .O(N__4653),
            .I(\Game_Inst.N_132 ));
    CascadeMux I__653 (
            .O(N__4646),
            .I(\Game_Inst.N_132_cascade_ ));
    InMux I__652 (
            .O(N__4643),
            .I(N__4639));
    InMux I__651 (
            .O(N__4642),
            .I(N__4636));
    LocalMux I__650 (
            .O(N__4639),
            .I(\Game_Inst.w_LFSR_Data_14 ));
    LocalMux I__649 (
            .O(N__4636),
            .I(\Game_Inst.w_LFSR_Data_14 ));
    CascadeMux I__648 (
            .O(N__4631),
            .I(N__4628));
    InMux I__647 (
            .O(N__4628),
            .I(N__4625));
    LocalMux I__646 (
            .O(N__4625),
            .I(N__4622));
    Odrv4 I__645 (
            .O(N__4622),
            .I(\Game_Inst.N_262 ));
    InMux I__644 (
            .O(N__4619),
            .I(N__4616));
    LocalMux I__643 (
            .O(N__4616),
            .I(N__4613));
    Odrv4 I__642 (
            .O(N__4613),
            .I(\Game_Inst.r_SM_Main_ns_i_i_a2_1_0_1 ));
    CascadeMux I__641 (
            .O(N__4610),
            .I(\Game_Inst.r_SM_Main_ns_i_i_1_1_cascade_ ));
    CascadeMux I__640 (
            .O(N__4607),
            .I(\Game_Inst.r_SM_Main_ns_i_i_3_1_cascade_ ));
    InMux I__639 (
            .O(N__4604),
            .I(N__4600));
    InMux I__638 (
            .O(N__4603),
            .I(N__4595));
    LocalMux I__637 (
            .O(N__4600),
            .I(N__4592));
    InMux I__636 (
            .O(N__4599),
            .I(N__4587));
    InMux I__635 (
            .O(N__4598),
            .I(N__4587));
    LocalMux I__634 (
            .O(N__4595),
            .I(\Game_Inst.N_137 ));
    Odrv4 I__633 (
            .O(N__4592),
            .I(\Game_Inst.N_137 ));
    LocalMux I__632 (
            .O(N__4587),
            .I(\Game_Inst.N_137 ));
    InMux I__631 (
            .O(N__4580),
            .I(N__4577));
    LocalMux I__630 (
            .O(N__4577),
            .I(N__4574));
    Odrv4 I__629 (
            .O(N__4574),
            .I(\Game_Inst.N_128 ));
    InMux I__628 (
            .O(N__4571),
            .I(N__4563));
    InMux I__627 (
            .O(N__4570),
            .I(N__4563));
    InMux I__626 (
            .O(N__4569),
            .I(N__4558));
    InMux I__625 (
            .O(N__4568),
            .I(N__4558));
    LocalMux I__624 (
            .O(N__4563),
            .I(\Game_Inst.N_91_2 ));
    LocalMux I__623 (
            .O(N__4558),
            .I(\Game_Inst.N_91_2 ));
    CascadeMux I__622 (
            .O(N__4553),
            .I(\Game_Inst.N_210_cascade_ ));
    InMux I__621 (
            .O(N__4550),
            .I(N__4544));
    InMux I__620 (
            .O(N__4549),
            .I(N__4544));
    LocalMux I__619 (
            .O(N__4544),
            .I(\Game_Inst.SUM_i_i_0_1 ));
    InMux I__618 (
            .O(N__4541),
            .I(N__4538));
    LocalMux I__617 (
            .O(N__4538),
            .I(N__4535));
    Odrv4 I__616 (
            .O(N__4535),
            .I(\Game_Inst.r_Pattern_0Z0Z_0 ));
    InMux I__615 (
            .O(N__4532),
            .I(N__4529));
    LocalMux I__614 (
            .O(N__4529),
            .I(\Game_Inst.r_Pattern_1Z0Z_0 ));
    CascadeMux I__613 (
            .O(N__4526),
            .I(\Game_Inst.r_Pattern_0_RNIDQ911Z0Z_0_cascade_ ));
    CascadeMux I__612 (
            .O(N__4523),
            .I(\Game_Inst.un6_r_button_dv_7_i_m2_ns_1_0_cascade_ ));
    InMux I__611 (
            .O(N__4520),
            .I(N__4517));
    LocalMux I__610 (
            .O(N__4517),
            .I(\Game_Inst.N_145 ));
    CascadeMux I__609 (
            .O(N__4514),
            .I(N__4511));
    InMux I__608 (
            .O(N__4511),
            .I(N__4508));
    LocalMux I__607 (
            .O(N__4508),
            .I(\Game_Inst.SUM_i_i_0_tz_0 ));
    InMux I__606 (
            .O(N__4505),
            .I(N__4500));
    InMux I__605 (
            .O(N__4504),
            .I(N__4495));
    InMux I__604 (
            .O(N__4503),
            .I(N__4495));
    LocalMux I__603 (
            .O(N__4500),
            .I(\Game_Inst.N_91 ));
    LocalMux I__602 (
            .O(N__4495),
            .I(\Game_Inst.N_91 ));
    CascadeMux I__601 (
            .O(N__4490),
            .I(\Game_Inst.r_SM_Main_ns_i_i_o2_0_1_1_cascade_ ));
    CascadeMux I__600 (
            .O(N__4487),
            .I(\Game_Inst.N_128_cascade_ ));
    InMux I__599 (
            .O(N__4484),
            .I(N__4478));
    InMux I__598 (
            .O(N__4483),
            .I(N__4478));
    LocalMux I__597 (
            .O(N__4478),
            .I(\Game_Inst.N_130 ));
    CascadeMux I__596 (
            .O(N__4475),
            .I(\Game_Inst.N_130_cascade_ ));
    InMux I__595 (
            .O(N__4472),
            .I(N__4469));
    LocalMux I__594 (
            .O(N__4469),
            .I(\Game_Inst.r_Index_0_sqmuxa_2_i_2_0 ));
    CascadeMux I__593 (
            .O(N__4466),
            .I(\Game_Inst.r_Index_0_sqmuxa_2_i_1_0_cascade_ ));
    CascadeMux I__592 (
            .O(N__4463),
            .I(\Game_Inst.N_209_cascade_ ));
    InMux I__591 (
            .O(N__4460),
            .I(N__4456));
    InMux I__590 (
            .O(N__4459),
            .I(N__4453));
    LocalMux I__589 (
            .O(N__4456),
            .I(N__4450));
    LocalMux I__588 (
            .O(N__4453),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_14 ));
    Odrv4 I__587 (
            .O(N__4450),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_14 ));
    InMux I__586 (
            .O(N__4445),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_13 ));
    InMux I__585 (
            .O(N__4442),
            .I(N__4438));
    InMux I__584 (
            .O(N__4441),
            .I(N__4435));
    LocalMux I__583 (
            .O(N__4438),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_15 ));
    LocalMux I__582 (
            .O(N__4435),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_15 ));
    InMux I__581 (
            .O(N__4430),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_14 ));
    InMux I__580 (
            .O(N__4427),
            .I(N__4423));
    InMux I__579 (
            .O(N__4426),
            .I(N__4420));
    LocalMux I__578 (
            .O(N__4423),
            .I(N__4417));
    LocalMux I__577 (
            .O(N__4420),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_16 ));
    Odrv4 I__576 (
            .O(N__4417),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_16 ));
    InMux I__575 (
            .O(N__4412),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_15 ));
    InMux I__574 (
            .O(N__4409),
            .I(N__4405));
    InMux I__573 (
            .O(N__4408),
            .I(N__4402));
    LocalMux I__572 (
            .O(N__4405),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_17 ));
    LocalMux I__571 (
            .O(N__4402),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_17 ));
    InMux I__570 (
            .O(N__4397),
            .I(bfn_6_8_0_));
    InMux I__569 (
            .O(N__4394),
            .I(N__4390));
    InMux I__568 (
            .O(N__4393),
            .I(N__4387));
    LocalMux I__567 (
            .O(N__4390),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_18 ));
    LocalMux I__566 (
            .O(N__4387),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_18 ));
    InMux I__565 (
            .O(N__4382),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_17 ));
    InMux I__564 (
            .O(N__4379),
            .I(N__4375));
    InMux I__563 (
            .O(N__4378),
            .I(N__4372));
    LocalMux I__562 (
            .O(N__4375),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_19 ));
    LocalMux I__561 (
            .O(N__4372),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_19 ));
    InMux I__560 (
            .O(N__4367),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_18 ));
    InMux I__559 (
            .O(N__4364),
            .I(N__4360));
    InMux I__558 (
            .O(N__4363),
            .I(N__4357));
    LocalMux I__557 (
            .O(N__4360),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_20 ));
    LocalMux I__556 (
            .O(N__4357),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_20 ));
    InMux I__555 (
            .O(N__4352),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_19 ));
    InMux I__554 (
            .O(N__4349),
            .I(N__4345));
    InMux I__553 (
            .O(N__4348),
            .I(N__4342));
    LocalMux I__552 (
            .O(N__4345),
            .I(N__4339));
    LocalMux I__551 (
            .O(N__4342),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_21 ));
    Odrv4 I__550 (
            .O(N__4339),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_21 ));
    InMux I__549 (
            .O(N__4334),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_20 ));
    InMux I__548 (
            .O(N__4331),
            .I(N__4310));
    InMux I__547 (
            .O(N__4330),
            .I(N__4310));
    InMux I__546 (
            .O(N__4329),
            .I(N__4310));
    InMux I__545 (
            .O(N__4328),
            .I(N__4310));
    InMux I__544 (
            .O(N__4327),
            .I(N__4307));
    InMux I__543 (
            .O(N__4326),
            .I(N__4302));
    InMux I__542 (
            .O(N__4325),
            .I(N__4302));
    InMux I__541 (
            .O(N__4324),
            .I(N__4299));
    InMux I__540 (
            .O(N__4323),
            .I(N__4294));
    InMux I__539 (
            .O(N__4322),
            .I(N__4294));
    InMux I__538 (
            .O(N__4321),
            .I(N__4287));
    InMux I__537 (
            .O(N__4320),
            .I(N__4287));
    InMux I__536 (
            .O(N__4319),
            .I(N__4287));
    LocalMux I__535 (
            .O(N__4310),
            .I(N__4282));
    LocalMux I__534 (
            .O(N__4307),
            .I(N__4282));
    LocalMux I__533 (
            .O(N__4302),
            .I(\Game_Inst.Count_Inst.un4_i_enable ));
    LocalMux I__532 (
            .O(N__4299),
            .I(\Game_Inst.Count_Inst.un4_i_enable ));
    LocalMux I__531 (
            .O(N__4294),
            .I(\Game_Inst.Count_Inst.un4_i_enable ));
    LocalMux I__530 (
            .O(N__4287),
            .I(\Game_Inst.Count_Inst.un4_i_enable ));
    Odrv4 I__529 (
            .O(N__4282),
            .I(\Game_Inst.Count_Inst.un4_i_enable ));
    InMux I__528 (
            .O(N__4271),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_21 ));
    CascadeMux I__527 (
            .O(N__4268),
            .I(N__4264));
    InMux I__526 (
            .O(N__4267),
            .I(N__4261));
    InMux I__525 (
            .O(N__4264),
            .I(N__4258));
    LocalMux I__524 (
            .O(N__4261),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_22 ));
    LocalMux I__523 (
            .O(N__4258),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_22 ));
    CEMux I__522 (
            .O(N__4253),
            .I(N__4241));
    CEMux I__521 (
            .O(N__4252),
            .I(N__4241));
    CEMux I__520 (
            .O(N__4251),
            .I(N__4241));
    CEMux I__519 (
            .O(N__4250),
            .I(N__4241));
    GlobalMux I__518 (
            .O(N__4241),
            .I(N__4238));
    gio2CtrlBuf I__517 (
            .O(N__4238),
            .I(\Game_Inst.N_83_i_g ));
    InMux I__516 (
            .O(N__4235),
            .I(N__4231));
    InMux I__515 (
            .O(N__4234),
            .I(N__4228));
    LocalMux I__514 (
            .O(N__4231),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_6 ));
    LocalMux I__513 (
            .O(N__4228),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_6 ));
    InMux I__512 (
            .O(N__4223),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_5 ));
    InMux I__511 (
            .O(N__4220),
            .I(N__4216));
    InMux I__510 (
            .O(N__4219),
            .I(N__4213));
    LocalMux I__509 (
            .O(N__4216),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_7 ));
    LocalMux I__508 (
            .O(N__4213),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_7 ));
    InMux I__507 (
            .O(N__4208),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_6 ));
    CascadeMux I__506 (
            .O(N__4205),
            .I(N__4201));
    InMux I__505 (
            .O(N__4204),
            .I(N__4198));
    InMux I__504 (
            .O(N__4201),
            .I(N__4195));
    LocalMux I__503 (
            .O(N__4198),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_8 ));
    LocalMux I__502 (
            .O(N__4195),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_8 ));
    InMux I__501 (
            .O(N__4190),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_7 ));
    InMux I__500 (
            .O(N__4187),
            .I(N__4183));
    InMux I__499 (
            .O(N__4186),
            .I(N__4180));
    LocalMux I__498 (
            .O(N__4183),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_9 ));
    LocalMux I__497 (
            .O(N__4180),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_9 ));
    InMux I__496 (
            .O(N__4175),
            .I(bfn_6_7_0_));
    InMux I__495 (
            .O(N__4172),
            .I(N__4168));
    InMux I__494 (
            .O(N__4171),
            .I(N__4165));
    LocalMux I__493 (
            .O(N__4168),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_10 ));
    LocalMux I__492 (
            .O(N__4165),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_10 ));
    InMux I__491 (
            .O(N__4160),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_9 ));
    InMux I__490 (
            .O(N__4157),
            .I(N__4153));
    InMux I__489 (
            .O(N__4156),
            .I(N__4150));
    LocalMux I__488 (
            .O(N__4153),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_11 ));
    LocalMux I__487 (
            .O(N__4150),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_11 ));
    InMux I__486 (
            .O(N__4145),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_10 ));
    CascadeMux I__485 (
            .O(N__4142),
            .I(N__4138));
    InMux I__484 (
            .O(N__4141),
            .I(N__4135));
    InMux I__483 (
            .O(N__4138),
            .I(N__4132));
    LocalMux I__482 (
            .O(N__4135),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_12 ));
    LocalMux I__481 (
            .O(N__4132),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_12 ));
    InMux I__480 (
            .O(N__4127),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_11 ));
    InMux I__479 (
            .O(N__4124),
            .I(N__4120));
    InMux I__478 (
            .O(N__4123),
            .I(N__4117));
    LocalMux I__477 (
            .O(N__4120),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_13 ));
    LocalMux I__476 (
            .O(N__4117),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_13 ));
    InMux I__475 (
            .O(N__4112),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_12 ));
    InMux I__474 (
            .O(N__4109),
            .I(N__4103));
    InMux I__473 (
            .O(N__4108),
            .I(N__4103));
    LocalMux I__472 (
            .O(N__4103),
            .I(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_20 ));
    InMux I__471 (
            .O(N__4100),
            .I(N__4097));
    LocalMux I__470 (
            .O(N__4097),
            .I(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_21 ));
    IoInMux I__469 (
            .O(N__4094),
            .I(N__4091));
    LocalMux I__468 (
            .O(N__4091),
            .I(N__4088));
    Odrv4 I__467 (
            .O(N__4088),
            .I(r_Hex_Encoding_i_2));
    InMux I__466 (
            .O(N__4085),
            .I(N__4080));
    InMux I__465 (
            .O(N__4084),
            .I(N__4077));
    InMux I__464 (
            .O(N__4083),
            .I(N__4074));
    LocalMux I__463 (
            .O(N__4080),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_1 ));
    LocalMux I__462 (
            .O(N__4077),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_1 ));
    LocalMux I__461 (
            .O(N__4074),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_1 ));
    CascadeMux I__460 (
            .O(N__4067),
            .I(N__4062));
    InMux I__459 (
            .O(N__4066),
            .I(N__4056));
    InMux I__458 (
            .O(N__4065),
            .I(N__4056));
    InMux I__457 (
            .O(N__4062),
            .I(N__4053));
    InMux I__456 (
            .O(N__4061),
            .I(N__4050));
    LocalMux I__455 (
            .O(N__4056),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_0 ));
    LocalMux I__454 (
            .O(N__4053),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_0 ));
    LocalMux I__453 (
            .O(N__4050),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_0 ));
    InMux I__452 (
            .O(N__4043),
            .I(N__4039));
    InMux I__451 (
            .O(N__4042),
            .I(N__4036));
    LocalMux I__450 (
            .O(N__4039),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_2 ));
    LocalMux I__449 (
            .O(N__4036),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_2 ));
    InMux I__448 (
            .O(N__4031),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_1 ));
    InMux I__447 (
            .O(N__4028),
            .I(N__4024));
    InMux I__446 (
            .O(N__4027),
            .I(N__4021));
    LocalMux I__445 (
            .O(N__4024),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_3 ));
    LocalMux I__444 (
            .O(N__4021),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_3 ));
    InMux I__443 (
            .O(N__4016),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_2 ));
    CascadeMux I__442 (
            .O(N__4013),
            .I(N__4010));
    InMux I__441 (
            .O(N__4010),
            .I(N__4006));
    InMux I__440 (
            .O(N__4009),
            .I(N__4003));
    LocalMux I__439 (
            .O(N__4006),
            .I(N__4000));
    LocalMux I__438 (
            .O(N__4003),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_4 ));
    Odrv4 I__437 (
            .O(N__4000),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_4 ));
    InMux I__436 (
            .O(N__3995),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_3 ));
    InMux I__435 (
            .O(N__3992),
            .I(N__3988));
    InMux I__434 (
            .O(N__3991),
            .I(N__3985));
    LocalMux I__433 (
            .O(N__3988),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_5 ));
    LocalMux I__432 (
            .O(N__3985),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_5 ));
    InMux I__431 (
            .O(N__3980),
            .I(\Game_Inst.Count_Inst.un2_r_counter_cry_4 ));
    InMux I__430 (
            .O(N__3977),
            .I(N__3974));
    LocalMux I__429 (
            .O(N__3974),
            .I(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_16 ));
    InMux I__428 (
            .O(N__3971),
            .I(N__3968));
    LocalMux I__427 (
            .O(N__3968),
            .I(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_17 ));
    InMux I__426 (
            .O(N__3965),
            .I(N__3962));
    LocalMux I__425 (
            .O(N__3962),
            .I(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_18 ));
    InMux I__424 (
            .O(N__3959),
            .I(N__3956));
    LocalMux I__423 (
            .O(N__3956),
            .I(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_19 ));
    InMux I__422 (
            .O(N__3953),
            .I(N__3950));
    LocalMux I__421 (
            .O(N__3950),
            .I(N__3946));
    InMux I__420 (
            .O(N__3949),
            .I(N__3943));
    Odrv4 I__419 (
            .O(N__3946),
            .I(\Game_Inst.w_LFSR_Data_0 ));
    LocalMux I__418 (
            .O(N__3943),
            .I(\Game_Inst.w_LFSR_Data_0 ));
    CascadeMux I__417 (
            .O(N__3938),
            .I(\Game_Inst.r_SM_Main_ns_i_0_a2_0_0_0_cascade_ ));
    InMux I__416 (
            .O(N__3935),
            .I(N__3932));
    LocalMux I__415 (
            .O(N__3932),
            .I(\Game_Inst.N_346 ));
    CascadeMux I__414 (
            .O(N__3929),
            .I(\Game_Inst.N_346_cascade_ ));
    CascadeMux I__413 (
            .O(N__3926),
            .I(N__3923));
    InMux I__412 (
            .O(N__3923),
            .I(N__3919));
    InMux I__411 (
            .O(N__3922),
            .I(N__3916));
    LocalMux I__410 (
            .O(N__3919),
            .I(\Game_Inst.o_Toggle_4_i_43 ));
    LocalMux I__409 (
            .O(N__3916),
            .I(\Game_Inst.o_Toggle_4_i_43 ));
    InMux I__408 (
            .O(N__3911),
            .I(N__3907));
    InMux I__407 (
            .O(N__3910),
            .I(N__3904));
    LocalMux I__406 (
            .O(N__3907),
            .I(\Debounce_SW1.r_CountZ0Z_6 ));
    LocalMux I__405 (
            .O(N__3904),
            .I(\Debounce_SW1.r_CountZ0Z_6 ));
    InMux I__404 (
            .O(N__3899),
            .I(N__3895));
    InMux I__403 (
            .O(N__3898),
            .I(N__3892));
    LocalMux I__402 (
            .O(N__3895),
            .I(\Debounce_SW1.r_CountZ0Z_5 ));
    LocalMux I__401 (
            .O(N__3892),
            .I(\Debounce_SW1.r_CountZ0Z_5 ));
    InMux I__400 (
            .O(N__3887),
            .I(N__3883));
    InMux I__399 (
            .O(N__3886),
            .I(N__3880));
    LocalMux I__398 (
            .O(N__3883),
            .I(\Debounce_SW1.r_CountZ0Z_4 ));
    LocalMux I__397 (
            .O(N__3880),
            .I(\Debounce_SW1.r_CountZ0Z_4 ));
    InMux I__396 (
            .O(N__3875),
            .I(N__3871));
    InMux I__395 (
            .O(N__3874),
            .I(N__3868));
    LocalMux I__394 (
            .O(N__3871),
            .I(\Debounce_SW1.r_CountZ0Z_16 ));
    LocalMux I__393 (
            .O(N__3868),
            .I(\Debounce_SW1.r_CountZ0Z_16 ));
    InMux I__392 (
            .O(N__3863),
            .I(N__3859));
    InMux I__391 (
            .O(N__3862),
            .I(N__3856));
    LocalMux I__390 (
            .O(N__3859),
            .I(\Debounce_SW1.r_CountZ0Z_15 ));
    LocalMux I__389 (
            .O(N__3856),
            .I(\Debounce_SW1.r_CountZ0Z_15 ));
    CascadeMux I__388 (
            .O(N__3851),
            .I(N__3848));
    InMux I__387 (
            .O(N__3848),
            .I(N__3844));
    InMux I__386 (
            .O(N__3847),
            .I(N__3841));
    LocalMux I__385 (
            .O(N__3844),
            .I(N__3838));
    LocalMux I__384 (
            .O(N__3841),
            .I(\Debounce_SW1.r_CountZ0Z_17 ));
    Odrv4 I__383 (
            .O(N__3838),
            .I(\Debounce_SW1.r_CountZ0Z_17 ));
    InMux I__382 (
            .O(N__3833),
            .I(N__3829));
    InMux I__381 (
            .O(N__3832),
            .I(N__3826));
    LocalMux I__380 (
            .O(N__3829),
            .I(\Debounce_SW1.r_CountZ0Z_14 ));
    LocalMux I__379 (
            .O(N__3826),
            .I(\Debounce_SW1.r_CountZ0Z_14 ));
    CascadeMux I__378 (
            .O(N__3821),
            .I(\Game_Inst.Count_Inst.un4_i_enable_16_cascade_ ));
    InMux I__377 (
            .O(N__3818),
            .I(N__3815));
    LocalMux I__376 (
            .O(N__3815),
            .I(\Game_Inst.Count_Inst.un4_i_enable_8 ));
    InMux I__375 (
            .O(N__3812),
            .I(N__3809));
    LocalMux I__374 (
            .O(N__3809),
            .I(\Game_Inst.Count_Inst.un4_i_enable_17 ));
    InMux I__373 (
            .O(N__3806),
            .I(N__3803));
    LocalMux I__372 (
            .O(N__3803),
            .I(N__3800));
    Odrv4 I__371 (
            .O(N__3800),
            .I(\Game_Inst.Count_Inst.un4_i_enable_14 ));
    CascadeMux I__370 (
            .O(N__3797),
            .I(\Game_Inst.Count_Inst.un4_i_enable_19_cascade_ ));
    InMux I__369 (
            .O(N__3794),
            .I(N__3791));
    LocalMux I__368 (
            .O(N__3791),
            .I(\Game_Inst.Count_Inst.un4_i_enable_13 ));
    InMux I__367 (
            .O(N__3788),
            .I(N__3784));
    InMux I__366 (
            .O(N__3787),
            .I(N__3781));
    LocalMux I__365 (
            .O(N__3784),
            .I(\Debounce_SW1.r_CountZ0Z_10 ));
    LocalMux I__364 (
            .O(N__3781),
            .I(\Debounce_SW1.r_CountZ0Z_10 ));
    InMux I__363 (
            .O(N__3776),
            .I(N__3772));
    InMux I__362 (
            .O(N__3775),
            .I(N__3769));
    LocalMux I__361 (
            .O(N__3772),
            .I(\Debounce_SW1.r_CountZ0Z_9 ));
    LocalMux I__360 (
            .O(N__3769),
            .I(\Debounce_SW1.r_CountZ0Z_9 ));
    CascadeMux I__359 (
            .O(N__3764),
            .I(N__3760));
    InMux I__358 (
            .O(N__3763),
            .I(N__3757));
    InMux I__357 (
            .O(N__3760),
            .I(N__3754));
    LocalMux I__356 (
            .O(N__3757),
            .I(\Debounce_SW1.r_CountZ0Z_11 ));
    LocalMux I__355 (
            .O(N__3754),
            .I(\Debounce_SW1.r_CountZ0Z_11 ));
    InMux I__354 (
            .O(N__3749),
            .I(N__3745));
    InMux I__353 (
            .O(N__3748),
            .I(N__3742));
    LocalMux I__352 (
            .O(N__3745),
            .I(\Debounce_SW1.r_CountZ0Z_8 ));
    LocalMux I__351 (
            .O(N__3742),
            .I(\Debounce_SW1.r_CountZ0Z_8 ));
    IoInMux I__350 (
            .O(N__3737),
            .I(N__3734));
    LocalMux I__349 (
            .O(N__3734),
            .I(r_Hex_Encoding_i_4));
    IoInMux I__348 (
            .O(N__3731),
            .I(N__3728));
    LocalMux I__347 (
            .O(N__3728),
            .I(N__3725));
    Span4Mux_s0_v I__346 (
            .O(N__3725),
            .I(N__3722));
    Odrv4 I__345 (
            .O(N__3722),
            .I(r_Hex_Encoding_i_5));
    IoInMux I__344 (
            .O(N__3719),
            .I(N__3716));
    LocalMux I__343 (
            .O(N__3716),
            .I(N__3713));
    Span4Mux_s0_v I__342 (
            .O(N__3713),
            .I(N__3710));
    Odrv4 I__341 (
            .O(N__3710),
            .I(r_Hex_Encoding_i_6));
    IoInMux I__340 (
            .O(N__3707),
            .I(N__3704));
    LocalMux I__339 (
            .O(N__3704),
            .I(r_Hex_Encoding_i_0));
    IoInMux I__338 (
            .O(N__3701),
            .I(N__3698));
    LocalMux I__337 (
            .O(N__3698),
            .I(r_Hex_Encoding_i_3));
    CascadeMux I__336 (
            .O(N__3695),
            .I(\Game_Inst.Count_Inst.un4_i_enable_12_cascade_ ));
    InMux I__335 (
            .O(N__3692),
            .I(\Debounce_SW1.un2_r_count_cry_10 ));
    InMux I__334 (
            .O(N__3689),
            .I(\Debounce_SW1.un2_r_count_cry_11 ));
    InMux I__333 (
            .O(N__3686),
            .I(\Debounce_SW1.un2_r_count_cry_12 ));
    InMux I__332 (
            .O(N__3683),
            .I(\Debounce_SW1.un2_r_count_cry_13 ));
    InMux I__331 (
            .O(N__3680),
            .I(\Debounce_SW1.un2_r_count_cry_14 ));
    InMux I__330 (
            .O(N__3677),
            .I(\Debounce_SW1.un2_r_count_cry_15 ));
    InMux I__329 (
            .O(N__3674),
            .I(bfn_4_9_0_));
    IoInMux I__328 (
            .O(N__3671),
            .I(N__3668));
    LocalMux I__327 (
            .O(N__3668),
            .I(N__3665));
    Span4Mux_s3_h I__326 (
            .O(N__3665),
            .I(N__3662));
    Odrv4 I__325 (
            .O(N__3662),
            .I(\Game_Inst.N_83_i ));
    IoInMux I__324 (
            .O(N__3659),
            .I(N__3656));
    LocalMux I__323 (
            .O(N__3656),
            .I(N__3653));
    Odrv12 I__322 (
            .O(N__3653),
            .I(r_Hex_Encoding_i_1));
    InMux I__321 (
            .O(N__3650),
            .I(\Debounce_SW1.un2_r_count_cry_1 ));
    InMux I__320 (
            .O(N__3647),
            .I(\Debounce_SW1.un2_r_count_cry_2 ));
    InMux I__319 (
            .O(N__3644),
            .I(\Debounce_SW1.un2_r_count_cry_3 ));
    InMux I__318 (
            .O(N__3641),
            .I(\Debounce_SW1.un2_r_count_cry_4 ));
    InMux I__317 (
            .O(N__3638),
            .I(\Debounce_SW1.un2_r_count_cry_5 ));
    InMux I__316 (
            .O(N__3635),
            .I(\Debounce_SW1.un2_r_count_cry_6 ));
    InMux I__315 (
            .O(N__3632),
            .I(\Debounce_SW1.un2_r_count_cry_7 ));
    InMux I__314 (
            .O(N__3629),
            .I(bfn_4_8_0_));
    InMux I__313 (
            .O(N__3626),
            .I(\Debounce_SW1.un2_r_count_cry_9 ));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(\Game_Inst.Count_Inst.un2_r_counter_cry_8 ),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_6_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_8_0_ (
            .carryinitin(\Game_Inst.Count_Inst.un2_r_counter_cry_16 ),
            .carryinitout(bfn_6_8_0_));
    defparam IN_MUX_bfv_7_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_5_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(\Debounce_SW4.un2_r_count_cry_8 ),
            .carryinitout(bfn_7_6_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(\Debounce_SW4.un2_r_count_cry_16 ),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(\Debounce_SW3.un2_r_count_cry_8 ),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(\Debounce_SW3.un2_r_count_cry_16 ),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\Debounce_SW2.un2_r_count_cry_8 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(\Debounce_SW2.un2_r_count_cry_16 ),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_4_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_7_0_));
    defparam IN_MUX_bfv_4_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_8_0_ (
            .carryinitin(\Debounce_SW1.un2_r_count_cry_8 ),
            .carryinitout(bfn_4_8_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(\Debounce_SW1.un2_r_count_cry_16 ),
            .carryinitout(bfn_4_9_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    ICE_GB \Debounce_SW3.r_State_e_0_RNI8LTG1_0  (
            .USERSIGNALTOGLOBALBUFFER(N__7865),
            .GLOBALBUFFEROUTPUT(\Debounce_SW3.N_40_g ));
    ICE_GB \Debounce_SW2.r_State_e_0_RNIKLK44_0  (
            .USERSIGNALTOGLOBALBUFFER(N__6272),
            .GLOBALBUFFEROUTPUT(\Debounce_SW2.N_38_g ));
    ICE_GB \Debounce_SW4.r_State_e_0_RNISK6T2_0  (
            .USERSIGNALTOGLOBALBUFFER(N__4778),
            .GLOBALBUFFEROUTPUT(\Debounce_SW4.N_42_g ));
    ICE_GB \Debounce_SW1.r_State_e_0_RNI0MBO2_0  (
            .USERSIGNALTOGLOBALBUFFER(N__5117),
            .GLOBALBUFFEROUTPUT(\Debounce_SW1.N_36_g ));
    GND GND (
            .Y(GNDG0));
    ICE_GB \Game_Inst.r_SM_Main_RNI9A2A_0_2  (
            .USERSIGNALTOGLOBALBUFFER(N__3671),
            .GLOBALBUFFEROUTPUT(\Game_Inst.N_83_i_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \Debounce_SW1.un2_r_count_cry_1_c_LC_4_7_0 .C_ON=1'b1;
    defparam \Debounce_SW1.un2_r_count_cry_1_c_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.un2_r_count_cry_1_c_LC_4_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Debounce_SW1.un2_r_count_cry_1_c_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(N__5879),
            .in2(N__5903),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_7_0_),
            .carryout(\Debounce_SW1.un2_r_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_2_LC_4_7_1 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_2_LC_4_7_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_2_LC_4_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_2_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(N__4945),
            .in2(_gnd_net_),
            .in3(N__3650),
            .lcout(\Debounce_SW1.r_CountZ0Z_2 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_1 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_2 ),
            .clk(N__8222),
            .ce(),
            .sr(N__5853));
    defparam \Debounce_SW1.r_Count_3_LC_4_7_2 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_3_LC_4_7_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_3_LC_4_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_3_LC_4_7_2  (
            .in0(_gnd_net_),
            .in1(N__4924),
            .in2(_gnd_net_),
            .in3(N__3647),
            .lcout(\Debounce_SW1.r_CountZ0Z_3 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_2 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_3 ),
            .clk(N__8222),
            .ce(),
            .sr(N__5853));
    defparam \Debounce_SW1.r_Count_4_LC_4_7_3 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_4_LC_4_7_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_4_LC_4_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_4_LC_4_7_3  (
            .in0(_gnd_net_),
            .in1(N__3887),
            .in2(_gnd_net_),
            .in3(N__3644),
            .lcout(\Debounce_SW1.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_3 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_4 ),
            .clk(N__8222),
            .ce(),
            .sr(N__5853));
    defparam \Debounce_SW1.r_Count_5_LC_4_7_4 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_5_LC_4_7_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_5_LC_4_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_5_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(N__3899),
            .in2(_gnd_net_),
            .in3(N__3641),
            .lcout(\Debounce_SW1.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_4 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_5 ),
            .clk(N__8222),
            .ce(),
            .sr(N__5853));
    defparam \Debounce_SW1.r_Count_6_LC_4_7_5 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_6_LC_4_7_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_6_LC_4_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_6_LC_4_7_5  (
            .in0(_gnd_net_),
            .in1(N__3911),
            .in2(_gnd_net_),
            .in3(N__3638),
            .lcout(\Debounce_SW1.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_5 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_6 ),
            .clk(N__8222),
            .ce(),
            .sr(N__5853));
    defparam \Debounce_SW1.r_Count_7_LC_4_7_6 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_7_LC_4_7_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_7_LC_4_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_7_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(N__5754),
            .in2(_gnd_net_),
            .in3(N__3635),
            .lcout(\Debounce_SW1.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_6 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_7 ),
            .clk(N__8222),
            .ce(),
            .sr(N__5853));
    defparam \Debounce_SW1.r_Count_8_LC_4_7_7 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_8_LC_4_7_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_8_LC_4_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_8_LC_4_7_7  (
            .in0(_gnd_net_),
            .in1(N__3749),
            .in2(_gnd_net_),
            .in3(N__3632),
            .lcout(\Debounce_SW1.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_7 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_8 ),
            .clk(N__8222),
            .ce(),
            .sr(N__5853));
    defparam \Debounce_SW1.r_Count_9_LC_4_8_0 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_9_LC_4_8_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_9_LC_4_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_9_LC_4_8_0  (
            .in0(_gnd_net_),
            .in1(N__3776),
            .in2(_gnd_net_),
            .in3(N__3629),
            .lcout(\Debounce_SW1.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_4_8_0_),
            .carryout(\Debounce_SW1.un2_r_count_cry_9 ),
            .clk(N__8221),
            .ce(),
            .sr(N__5852));
    defparam \Debounce_SW1.r_Count_10_LC_4_8_1 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_10_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_10_LC_4_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_10_LC_4_8_1  (
            .in0(_gnd_net_),
            .in1(N__3788),
            .in2(_gnd_net_),
            .in3(N__3626),
            .lcout(\Debounce_SW1.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_9 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_10 ),
            .clk(N__8221),
            .ce(),
            .sr(N__5852));
    defparam \Debounce_SW1.r_Count_11_LC_4_8_2 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_11_LC_4_8_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_11_LC_4_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_11_LC_4_8_2  (
            .in0(_gnd_net_),
            .in1(N__3763),
            .in2(_gnd_net_),
            .in3(N__3692),
            .lcout(\Debounce_SW1.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_10 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_11 ),
            .clk(N__8221),
            .ce(),
            .sr(N__5852));
    defparam \Debounce_SW1.r_Count_12_LC_4_8_3 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_12_LC_4_8_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_12_LC_4_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_12_LC_4_8_3  (
            .in0(_gnd_net_),
            .in1(N__5811),
            .in2(_gnd_net_),
            .in3(N__3689),
            .lcout(\Debounce_SW1.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_11 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_12 ),
            .clk(N__8221),
            .ce(),
            .sr(N__5852));
    defparam \Debounce_SW1.r_Count_13_LC_4_8_4 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_13_LC_4_8_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_13_LC_4_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_13_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(N__5781),
            .in2(_gnd_net_),
            .in3(N__3686),
            .lcout(\Debounce_SW1.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_12 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_13 ),
            .clk(N__8221),
            .ce(),
            .sr(N__5852));
    defparam \Debounce_SW1.r_Count_14_LC_4_8_5 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_14_LC_4_8_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_14_LC_4_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_14_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(N__3833),
            .in2(_gnd_net_),
            .in3(N__3683),
            .lcout(\Debounce_SW1.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_13 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_14 ),
            .clk(N__8221),
            .ce(),
            .sr(N__5852));
    defparam \Debounce_SW1.r_Count_15_LC_4_8_6 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_15_LC_4_8_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_15_LC_4_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_15_LC_4_8_6  (
            .in0(_gnd_net_),
            .in1(N__3863),
            .in2(_gnd_net_),
            .in3(N__3680),
            .lcout(\Debounce_SW1.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_14 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_15 ),
            .clk(N__8221),
            .ce(),
            .sr(N__5852));
    defparam \Debounce_SW1.r_Count_16_LC_4_8_7 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_16_LC_4_8_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_16_LC_4_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_16_LC_4_8_7  (
            .in0(_gnd_net_),
            .in1(N__3875),
            .in2(_gnd_net_),
            .in3(N__3677),
            .lcout(\Debounce_SW1.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Debounce_SW1.un2_r_count_cry_15 ),
            .carryout(\Debounce_SW1.un2_r_count_cry_16 ),
            .clk(N__8221),
            .ce(),
            .sr(N__5852));
    defparam \Debounce_SW1.r_Count_17_LC_4_9_0 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_17_LC_4_9_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_17_LC_4_9_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Debounce_SW1.r_Count_17_LC_4_9_0  (
            .in0(_gnd_net_),
            .in1(N__3847),
            .in2(_gnd_net_),
            .in3(N__3674),
            .lcout(\Debounce_SW1.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8223),
            .ce(),
            .sr(N__5854));
    defparam \Game_Inst.r_SM_Main_RNI9A2A_2_LC_4_10_5 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI9A2A_2_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI9A2A_2_LC_4_10_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Game_Inst.r_SM_Main_RNI9A2A_2_LC_4_10_5  (
            .in0(_gnd_net_),
            .in1(N__3922),
            .in2(_gnd_net_),
            .in3(N__7603),
            .lcout(\Game_Inst.N_83_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_1_LC_4_12_0 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_1_LC_4_12_0 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_1_LC_4_12_0 .LUT_INIT=16'b0010110100000100;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_1_LC_4_12_0  (
            .in0(N__7235),
            .in1(N__7830),
            .in2(N__6956),
            .in3(N__7761),
            .lcout(r_Hex_Encoding_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8230),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_4_LC_4_16_0 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_4_LC_4_16_0 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_4_LC_4_16_0 .LUT_INIT=16'b1100010000010000;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_4_LC_4_16_0  (
            .in0(N__7764),
            .in1(N__7251),
            .in2(N__7852),
            .in3(N__6967),
            .lcout(r_Hex_Encoding_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8254),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_5_LC_4_16_1 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_5_LC_4_16_1 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_5_LC_4_16_1 .LUT_INIT=16'b1100001010101000;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_5_LC_4_16_1  (
            .in0(N__7252),
            .in1(N__7845),
            .in2(N__6971),
            .in3(N__7765),
            .lcout(r_Hex_Encoding_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8254),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_6_LC_4_16_2 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_6_LC_4_16_2 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_6_LC_4_16_2 .LUT_INIT=16'b0010100000000110;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_6_LC_4_16_2  (
            .in0(N__7766),
            .in1(N__7253),
            .in2(N__7853),
            .in3(N__6968),
            .lcout(r_Hex_Encoding_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8254),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_0_LC_4_16_3 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_0_LC_4_16_3 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_0_LC_4_16_3 .LUT_INIT=16'b0000100100100001;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_0_LC_4_16_3  (
            .in0(N__7249),
            .in1(N__7843),
            .in2(N__6969),
            .in3(N__7762),
            .lcout(r_Hex_Encoding_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8254),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_3_LC_4_16_7 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_3_LC_4_16_7 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_3_LC_4_16_7 .LUT_INIT=16'b1000100101000010;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_3_LC_4_16_7  (
            .in0(N__7250),
            .in1(N__7844),
            .in2(N__6970),
            .in3(N__7763),
            .lcout(r_Hex_Encoding_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8254),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_0_LC_5_6_3 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_0_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_0_LC_5_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_0_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4065),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8227),
            .ce(N__4251),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_1_LC_5_6_7 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_1_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_1_LC_5_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_1_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(N__4066),
            .in2(_gnd_net_),
            .in3(N__4085),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8227),
            .ce(N__4251),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNI2H0N1_5_LC_5_7_0 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNI2H0N1_5_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNI2H0N1_5_LC_5_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNI2H0N1_5_LC_5_7_0  (
            .in0(N__4234),
            .in1(N__4219),
            .in2(N__4205),
            .in3(N__3991),
            .lcout(),
            .ltout(\Game_Inst.Count_Inst.un4_i_enable_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNI233G2_13_LC_5_7_1 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNI233G2_13_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNI233G2_13_LC_5_7_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNI233G2_13_LC_5_7_1  (
            .in0(N__4061),
            .in1(N__4441),
            .in2(N__3695),
            .in3(N__4123),
            .lcout(\Game_Inst.Count_Inst.un4_i_enable_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNII00N1_1_LC_5_7_3 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNII00N1_1_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNII00N1_1_LC_5_7_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNII00N1_1_LC_5_7_3  (
            .in0(N__4083),
            .in1(N__4027),
            .in2(N__4013),
            .in3(N__4042),
            .lcout(\Game_Inst.Count_Inst.un4_i_enable_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_RNIS1S7_4_LC_5_7_5 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_RNIS1S7_4_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_RNIS1S7_4_LC_5_7_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Debounce_SW1.r_Count_RNIS1S7_4_LC_5_7_5  (
            .in0(N__3910),
            .in1(N__3898),
            .in2(_gnd_net_),
            .in3(N__3886),
            .lcout(\Debounce_SW1.N_146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNI7SNU_10_LC_5_7_6 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNI7SNU_10_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNI7SNU_10_LC_5_7_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNI7SNU_10_LC_5_7_6  (
            .in0(N__4156),
            .in1(N__4171),
            .in2(N__4142),
            .in3(N__4186),
            .lcout(\Game_Inst.Count_Inst.un4_i_enable_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_RNIMQSP_17_LC_5_8_0 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_RNIMQSP_17_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_RNIMQSP_17_LC_5_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW1.r_Count_RNIMQSP_17_LC_5_8_0  (
            .in0(N__3874),
            .in1(N__3862),
            .in2(N__3851),
            .in3(N__3832),
            .lcout(\Debounce_SW1.r_count15_i_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNILRAB_17_LC_5_8_1 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNILRAB_17_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNILRAB_17_LC_5_8_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNILRAB_17_LC_5_8_1  (
            .in0(N__4393),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4408),
            .lcout(\Game_Inst.Count_Inst.un4_i_enable_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNIRAOM_22_LC_5_8_2 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIRAOM_22_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIRAOM_22_LC_5_8_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNIRAOM_22_LC_5_8_2  (
            .in0(N__4349),
            .in1(N__4363),
            .in2(N__4268),
            .in3(N__4378),
            .lcout(),
            .ltout(\Game_Inst.Count_Inst.un4_i_enable_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNI0TDD1_14_LC_5_8_3 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNI0TDD1_14_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNI0TDD1_14_LC_5_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNI0TDD1_14_LC_5_8_3  (
            .in0(N__4460),
            .in1(N__4427),
            .in2(N__3821),
            .in3(N__3818),
            .lcout(),
            .ltout(\Game_Inst.Count_Inst.un4_i_enable_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNIRS8J6_10_LC_5_8_4 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIRS8J6_10_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIRS8J6_10_LC_5_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNIRS8J6_10_LC_5_8_4  (
            .in0(N__3812),
            .in1(N__3806),
            .in2(N__3797),
            .in3(N__3794),
            .lcout(\Game_Inst.Count_Inst.un4_i_enable ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_RNIGB6I_8_LC_5_8_7 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_RNIGB6I_8_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_RNIGB6I_8_LC_5_8_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Debounce_SW1.r_Count_RNIGB6I_8_LC_5_8_7  (
            .in0(N__3787),
            .in1(N__3775),
            .in2(N__3764),
            .in3(N__3748),
            .lcout(\Debounce_SW1.N_161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.o_Toggle_LC_5_9_7 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.o_Toggle_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.o_Toggle_LC_5_9_7 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \Game_Inst.Count_Inst.o_Toggle_LC_5_9_7  (
            .in0(N__5643),
            .in1(N__7604),
            .in2(N__3926),
            .in3(N__4324),
            .lcout(\Game_Inst.w_Toggle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8225),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNO_0_0_LC_5_10_0 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNO_0_0_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNO_0_0_LC_5_10_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Game_Inst.r_Index_RNO_0_0_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__5166),
            .in2(_gnd_net_),
            .in3(N__3935),
            .lcout(\Game_Inst.SUM_i_i_0_tz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_1_0_LC_5_10_2 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_1_0_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_1_0_LC_5_10_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_1_0_LC_5_10_2  (
            .in0(N__7659),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4664),
            .lcout(),
            .ltout(\Game_Inst.r_SM_Main_ns_i_0_a2_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_0_LC_5_10_3 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_0_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_SM_Main_0_LC_5_10_3 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \Game_Inst.r_SM_Main_0_LC_5_10_3  (
            .in0(N__4484),
            .in1(N__4603),
            .in2(N__3938),
            .in3(N__5153),
            .lcout(\Game_Inst.r_SM_MainZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8226),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNIGERD7_0_LC_5_10_4 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNIGERD7_0_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNIGERD7_0_LC_5_10_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Game_Inst.r_SM_Main_RNIGERD7_0_LC_5_10_4  (
            .in0(N__7658),
            .in1(N__7479),
            .in2(N__7416),
            .in3(N__4483),
            .lcout(\Game_Inst.N_346 ),
            .ltout(\Game_Inst.N_346_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNICF6P8_1_LC_5_10_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNICF6P8_1_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNICF6P8_1_LC_5_10_5 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \Game_Inst.r_Index_RNICF6P8_1_LC_5_10_5  (
            .in0(N__5167),
            .in1(N__5249),
            .in2(N__3929),
            .in3(N__5339),
            .lcout(\Game_Inst.SUM_i_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.counter_o_Toggle_4_i_43_LC_5_10_7 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.counter_o_Toggle_4_i_43_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.counter_o_Toggle_4_i_43_LC_5_10_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \Game_Inst.Count_Inst.counter_o_Toggle_4_i_43_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(N__7398),
            .in2(_gnd_net_),
            .in3(N__7657),
            .lcout(\Game_Inst.o_Toggle_4_i_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_6_0_LC_5_11_0 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_6_0_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_6_0_LC_5_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_6_0_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7028),
            .lcout(\Game_Inst.r_Pattern_6Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8231),
            .ce(N__6067),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_0_0_LC_5_11_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_0_0_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_0_0_LC_5_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_0_0_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3953),
            .lcout(\Game_Inst.r_Pattern_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8231),
            .ce(N__6067),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_7_0_LC_5_11_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_7_0_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_7_0_LC_5_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_7_0_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4642),
            .lcout(\Game_Inst.r_Pattern_7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8231),
            .ce(N__6067),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_1_0_LC_5_11_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_1_0_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_1_0_LC_5_11_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \Game_Inst.r_Pattern_1_0_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__6014),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Game_Inst.r_Pattern_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8231),
            .ce(N__6067),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_1_LC_5_12_1 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_1_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_1_LC_5_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_1_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3949),
            .lcout(\Game_Inst.w_LFSR_Data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8237),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_16_LC_5_12_2 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_16_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_16_LC_5_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_16_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6097),
            .lcout(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8237),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_15_LC_5_12_3 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_15_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_15_LC_5_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_15_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4643),
            .lcout(\Game_Inst.w_LFSR_Data_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8237),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_20_LC_5_13_0 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_20_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_20_LC_5_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_20_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3959),
            .lcout(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8242),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_17_LC_5_13_1 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_17_LC_5_13_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_17_LC_5_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_17_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3977),
            .lcout(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8242),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_18_LC_5_13_2 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_18_LC_5_13_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_18_LC_5_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_18_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3971),
            .lcout(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8242),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_19_LC_5_13_5 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_19_LC_5_13_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_19_LC_5_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_19_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3965),
            .lcout(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8242),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_0_LC_5_13_6 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_0_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_0_LC_5_13_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_0_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(N__4100),
            .in2(_gnd_net_),
            .in3(N__4108),
            .lcout(\Game_Inst.w_LFSR_Data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8242),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_21_LC_5_13_7 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_21_LC_5_13_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_21_LC_5_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_21_LC_5_13_7  (
            .in0(N__4109),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8242),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_2_LC_5_15_5 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_2_LC_5_15_5 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_2_LC_5_15_5 .LUT_INIT=16'b0001111100000010;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_2_LC_5_15_5  (
            .in0(N__7237),
            .in1(N__7831),
            .in2(N__6957),
            .in3(N__7746),
            .lcout(r_Hex_Encoding_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8255),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_0_LC_6_4_0 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_0_LC_6_4_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_0_LC_6_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Debounce_SW4.r_Count_0_LC_6_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4732),
            .lcout(\Debounce_SW4.r_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8244),
            .ce(),
            .sr(N__4965));
    defparam \Debounce_SW4.r_Count_1_LC_6_4_1 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_1_LC_6_4_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_1_LC_6_4_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Debounce_SW4.r_Count_1_LC_6_4_1  (
            .in0(N__4733),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4711),
            .lcout(\Debounce_SW4.r_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8244),
            .ce(),
            .sr(N__4965));
    defparam \Game_Inst.Count_Inst.un2_r_counter_cry_1_c_LC_6_6_0 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.un2_r_counter_cry_1_c_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.un2_r_counter_cry_1_c_LC_6_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Game_Inst.Count_Inst.un2_r_counter_cry_1_c_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__4084),
            .in2(N__4067),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_2_LC_6_6_1 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_2_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_2_LC_6_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_2_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__4043),
            .in2(_gnd_net_),
            .in3(N__4031),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_2 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_1 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_2 ),
            .clk(N__8233),
            .ce(N__4253),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_3_LC_6_6_2 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_3_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_3_LC_6_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_3_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__4028),
            .in2(_gnd_net_),
            .in3(N__4016),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_3 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_2 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_3 ),
            .clk(N__8233),
            .ce(N__4253),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_4_LC_6_6_3 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_4_LC_6_6_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_4_LC_6_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_4_LC_6_6_3  (
            .in0(N__4327),
            .in1(N__4009),
            .in2(_gnd_net_),
            .in3(N__3995),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_4 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_3 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_4 ),
            .clk(N__8233),
            .ce(N__4253),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_5_LC_6_6_4 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_5_LC_6_6_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_5_LC_6_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_5_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(N__3992),
            .in2(_gnd_net_),
            .in3(N__3980),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_5 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_4 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_5 ),
            .clk(N__8233),
            .ce(N__4253),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_6_LC_6_6_5 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_6_LC_6_6_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_6_LC_6_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_6_LC_6_6_5  (
            .in0(_gnd_net_),
            .in1(N__4235),
            .in2(_gnd_net_),
            .in3(N__4223),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_6 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_5 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_6 ),
            .clk(N__8233),
            .ce(N__4253),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_7_LC_6_6_6 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_7_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_7_LC_6_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_7_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(N__4220),
            .in2(_gnd_net_),
            .in3(N__4208),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_7 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_6 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_7 ),
            .clk(N__8233),
            .ce(N__4253),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_8_LC_6_6_7 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_8_LC_6_6_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_8_LC_6_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_8_LC_6_6_7  (
            .in0(_gnd_net_),
            .in1(N__4204),
            .in2(_gnd_net_),
            .in3(N__4190),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_8 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_7 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_8 ),
            .clk(N__8233),
            .ce(N__4253),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_9_LC_6_7_0 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_9_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_9_LC_6_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_9_LC_6_7_0  (
            .in0(N__4323),
            .in1(N__4187),
            .in2(_gnd_net_),
            .in3(N__4175),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_9 ),
            .clk(N__8228),
            .ce(N__4252),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_10_LC_6_7_1 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_10_LC_6_7_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_10_LC_6_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_10_LC_6_7_1  (
            .in0(N__4328),
            .in1(N__4172),
            .in2(_gnd_net_),
            .in3(N__4160),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_10 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_9 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_10 ),
            .clk(N__8228),
            .ce(N__4252),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_11_LC_6_7_2 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_11_LC_6_7_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_11_LC_6_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_11_LC_6_7_2  (
            .in0(N__4322),
            .in1(N__4157),
            .in2(_gnd_net_),
            .in3(N__4145),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_11 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_10 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_11 ),
            .clk(N__8228),
            .ce(N__4252),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_12_LC_6_7_3 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_12_LC_6_7_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_12_LC_6_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_12_LC_6_7_3  (
            .in0(N__4329),
            .in1(N__4141),
            .in2(_gnd_net_),
            .in3(N__4127),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_12 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_11 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_12 ),
            .clk(N__8228),
            .ce(N__4252),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_13_LC_6_7_4 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_13_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_13_LC_6_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_13_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(N__4124),
            .in2(_gnd_net_),
            .in3(N__4112),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_13 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_12 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_13 ),
            .clk(N__8228),
            .ce(N__4252),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_14_LC_6_7_5 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_14_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_14_LC_6_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_14_LC_6_7_5  (
            .in0(N__4330),
            .in1(N__4459),
            .in2(_gnd_net_),
            .in3(N__4445),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_14 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_13 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_14 ),
            .clk(N__8228),
            .ce(N__4252),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_15_LC_6_7_6 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_15_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_15_LC_6_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_15_LC_6_7_6  (
            .in0(_gnd_net_),
            .in1(N__4442),
            .in2(_gnd_net_),
            .in3(N__4430),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_15 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_14 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_15 ),
            .clk(N__8228),
            .ce(N__4252),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_16_LC_6_7_7 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_16_LC_6_7_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_16_LC_6_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_16_LC_6_7_7  (
            .in0(N__4331),
            .in1(N__4426),
            .in2(_gnd_net_),
            .in3(N__4412),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_16 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_15 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_16 ),
            .clk(N__8228),
            .ce(N__4252),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_17_LC_6_8_0 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_17_LC_6_8_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_17_LC_6_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_17_LC_6_8_0  (
            .in0(N__4325),
            .in1(N__4409),
            .in2(_gnd_net_),
            .in3(N__4397),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_6_8_0_),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_17 ),
            .clk(N__8224),
            .ce(N__4250),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_18_LC_6_8_1 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_18_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_18_LC_6_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_18_LC_6_8_1  (
            .in0(N__4319),
            .in1(N__4394),
            .in2(_gnd_net_),
            .in3(N__4382),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_18 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_17 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_18 ),
            .clk(N__8224),
            .ce(N__4250),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_19_LC_6_8_2 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_19_LC_6_8_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_19_LC_6_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_19_LC_6_8_2  (
            .in0(N__4326),
            .in1(N__4379),
            .in2(_gnd_net_),
            .in3(N__4367),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_19 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_18 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_19 ),
            .clk(N__8224),
            .ce(N__4250),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_20_LC_6_8_3 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_20_LC_6_8_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_20_LC_6_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_20_LC_6_8_3  (
            .in0(N__4320),
            .in1(N__4364),
            .in2(_gnd_net_),
            .in3(N__4352),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_20 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_19 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_20 ),
            .clk(N__8224),
            .ce(N__4250),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_21_LC_6_8_4 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_21_LC_6_8_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_21_LC_6_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_21_LC_6_8_4  (
            .in0(_gnd_net_),
            .in1(N__4348),
            .in2(_gnd_net_),
            .in3(N__4334),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_21 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un2_r_counter_cry_20 ),
            .carryout(\Game_Inst.Count_Inst.un2_r_counter_cry_21 ),
            .clk(N__8224),
            .ce(N__4250),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_22_LC_6_8_5 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_22_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_22_LC_6_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_22_LC_6_8_5  (
            .in0(N__4321),
            .in1(N__4267),
            .in2(_gnd_net_),
            .in3(N__4271),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8224),
            .ce(N__4250),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNO_1_0_LC_6_9_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNO_1_0_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNO_1_0_LC_6_9_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Game_Inst.r_Index_RNO_1_0_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__4670),
            .in2(_gnd_net_),
            .in3(N__4569),
            .lcout(\Game_Inst.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_ID_RNIRM4R6_0_LC_6_9_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_ID_RNIRM4R6_0_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Button_ID_RNIRM4R6_0_LC_6_9_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Game_Inst.r_Button_ID_RNIRM4R6_0_LC_6_9_2  (
            .in0(N__5075),
            .in1(N__5108),
            .in2(N__8101),
            .in3(N__7960),
            .lcout(\Game_Inst.N_128 ),
            .ltout(\Game_Inst.N_128_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_DV_RNI62R37_LC_6_9_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_DV_RNI62R37_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Button_DV_RNI62R37_LC_6_9_3 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \Game_Inst.r_Button_DV_RNI62R37_LC_6_9_3  (
            .in0(N__5363),
            .in1(_gnd_net_),
            .in2(N__4487),
            .in3(_gnd_net_),
            .lcout(\Game_Inst.N_130 ),
            .ltout(\Game_Inst.N_130_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNIIOU38_0_LC_6_9_4 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNIIOU38_0_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNIIOU38_0_LC_6_9_4 .LUT_INIT=16'b1111110111101100;
    LogicCell40 \Game_Inst.r_SM_Main_RNIIOU38_0_LC_6_9_4  (
            .in0(N__7653),
            .in1(N__4472),
            .in2(N__4475),
            .in3(N__7602),
            .lcout(\Game_Inst.N_91_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Toggle_RNI6QCP_LC_6_9_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Toggle_RNI6QCP_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Toggle_RNI6QCP_LC_6_9_5 .LUT_INIT=16'b0011001111000100;
    LogicCell40 \Game_Inst.r_Toggle_RNI6QCP_LC_6_9_5  (
            .in0(N__5593),
            .in1(N__7402),
            .in2(N__5648),
            .in3(N__7652),
            .lcout(\Game_Inst.r_Index_0_sqmuxa_2_i_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_DV_RNIJABF_LC_6_9_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_DV_RNIJABF_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Button_DV_RNIJABF_LC_6_9_6 .LUT_INIT=16'b0000101010101110;
    LogicCell40 \Game_Inst.r_Button_DV_RNIJABF_LC_6_9_6  (
            .in0(N__7403),
            .in1(N__5364),
            .in2(N__8056),
            .in3(N__7114),
            .lcout(),
            .ltout(\Game_Inst.r_Index_0_sqmuxa_2_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNIRLCOA_1_LC_6_9_7 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNIRLCOA_1_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNIRLCOA_1_LC_6_9_7 .LUT_INIT=16'b1111111110001111;
    LogicCell40 \Game_Inst.r_SM_Main_RNIRLCOA_1_LC_6_9_7  (
            .in0(N__4604),
            .in1(N__7404),
            .in2(N__4466),
            .in3(N__4568),
            .lcout(\Game_Inst.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNO_0_1_LC_6_10_0 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNO_0_1_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNO_0_1_LC_6_10_0 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \Game_Inst.r_Index_RNO_0_1_LC_6_10_0  (
            .in0(N__5340),
            .in1(N__4668),
            .in2(_gnd_net_),
            .in3(N__4570),
            .lcout(),
            .ltout(\Game_Inst.N_209_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_1_LC_6_10_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_1_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Index_1_LC_6_10_1 .LUT_INIT=16'b0000000010001010;
    LogicCell40 \Game_Inst.r_Index_1_LC_6_10_1  (
            .in0(N__4505),
            .in1(N__5247),
            .in2(N__4463),
            .in3(N__4549),
            .lcout(\Game_Inst.r_IndexZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8232),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNO_0_2_LC_6_10_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNO_0_2_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNO_0_2_LC_6_10_2 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \Game_Inst.r_Index_RNO_0_2_LC_6_10_2  (
            .in0(N__5246),
            .in1(N__4669),
            .in2(N__5345),
            .in3(N__4571),
            .lcout(),
            .ltout(\Game_Inst.N_210_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_2_LC_6_10_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_2_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Index_2_LC_6_10_3 .LUT_INIT=16'b0000010010001100;
    LogicCell40 \Game_Inst.r_Index_2_LC_6_10_3  (
            .in0(N__5215),
            .in1(N__4504),
            .in2(N__4553),
            .in3(N__4550),
            .lcout(\Game_Inst.r_IndexZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8232),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_0_RNIDQ911_0_LC_6_10_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_0_RNIDQ911_0_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_0_RNIDQ911_0_LC_6_10_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Game_Inst.r_Pattern_0_RNIDQ911_0_LC_6_10_4  (
            .in0(N__4541),
            .in1(N__5338),
            .in2(_gnd_net_),
            .in3(N__4532),
            .lcout(),
            .ltout(\Game_Inst.r_Pattern_0_RNIDQ911Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNID9922_1_LC_6_10_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNID9922_1_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNID9922_1_LC_6_10_5 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \Game_Inst.r_Index_RNID9922_1_LC_6_10_5  (
            .in0(N__5213),
            .in1(N__5245),
            .in2(N__4526),
            .in3(N__5186),
            .lcout(),
            .ltout(\Game_Inst.un6_r_button_dv_7_i_m2_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNIJFF03_2_LC_6_10_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNIJFF03_2_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNIJFF03_2_LC_6_10_6 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \Game_Inst.r_Index_RNIJFF03_2_LC_6_10_6  (
            .in0(N__5282),
            .in1(N__4679),
            .in2(N__4523),
            .in3(N__5214),
            .lcout(\Game_Inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_0_LC_6_10_7 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_0_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Index_0_LC_6_10_7 .LUT_INIT=16'b0001110100000000;
    LogicCell40 \Game_Inst.r_Index_0_LC_6_10_7  (
            .in0(N__4520),
            .in1(N__5344),
            .in2(N__4514),
            .in3(N__4503),
            .lcout(\Game_Inst.r_IndexZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8232),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_4_1_LC_6_11_0 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_4_1_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_4_1_LC_6_11_0 .LUT_INIT=16'b0011000100000000;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_4_1_LC_6_11_0  (
            .in0(N__5601),
            .in1(N__7406),
            .in2(N__5665),
            .in3(N__7654),
            .lcout(\Game_Inst.N_262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNI2PL31_1_LC_6_11_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNI2PL31_1_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNI2PL31_1_LC_6_11_1 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \Game_Inst.r_Index_RNI2PL31_1_LC_6_11_1  (
            .in0(N__5332),
            .in1(N__7736),
            .in2(N__7829),
            .in3(N__5248),
            .lcout(),
            .ltout(\Game_Inst.r_SM_Main_ns_i_i_o2_0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNIJ4N12_2_LC_6_11_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNIJ4N12_2_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNIJ4N12_2_LC_6_11_2 .LUT_INIT=16'b1111101111111110;
    LogicCell40 \Game_Inst.r_Index_RNIJ4N12_2_LC_6_11_2  (
            .in0(N__6928),
            .in1(N__7236),
            .in2(N__4490),
            .in3(N__5216),
            .lcout(\Game_Inst.N_137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_2_1_LC_6_11_3 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_2_1_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_2_1_LC_6_11_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_2_1_LC_6_11_3  (
            .in0(N__7656),
            .in1(N__5603),
            .in2(N__5666),
            .in3(N__7559),
            .lcout(\Game_Inst.r_SM_Main_ns_i_i_a2_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_6_RNIPUEE_0_LC_6_11_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_6_RNIPUEE_0_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_6_RNIPUEE_0_LC_6_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Game_Inst.r_Pattern_6_RNIPUEE_0_LC_6_11_4  (
            .in0(N__4691),
            .in1(N__4685),
            .in2(_gnd_net_),
            .in3(N__5331),
            .lcout(\Game_Inst.r_Pattern_6_RNIPUEEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNICE0A_1_LC_6_11_5 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNICE0A_1_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNICE0A_1_LC_6_11_5 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \Game_Inst.r_SM_Main_RNICE0A_1_LC_6_11_5  (
            .in0(N__7405),
            .in1(N__8046),
            .in2(N__7583),
            .in3(N__7112),
            .lcout(\Game_Inst.N_132 ),
            .ltout(\Game_Inst.N_132_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Toggle_RNIFQ101_LC_6_11_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Toggle_RNIFQ101_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Toggle_RNIFQ101_LC_6_11_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Game_Inst.r_Toggle_RNIFQ101_LC_6_11_6  (
            .in0(N__5602),
            .in1(N__5661),
            .in2(N__4646),
            .in3(N__7655),
            .lcout(\Game_Inst.N_303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_14_LC_6_11_7 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_14_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_14_LC_6_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_14_LC_6_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7010),
            .lcout(\Game_Inst.w_LFSR_Data_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8238),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_1_1_LC_6_12_1 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_1_1_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_1_1_LC_6_12_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_1_1_LC_6_12_1  (
            .in0(N__7558),
            .in1(N__7484),
            .in2(N__4631),
            .in3(N__7679),
            .lcout(),
            .ltout(\Game_Inst.r_SM_Main_ns_i_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_0_1_LC_6_12_2 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_0_1_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_0_1_LC_6_12_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_0_1_LC_6_12_2  (
            .in0(N__4599),
            .in1(N__4619),
            .in2(N__4610),
            .in3(N__5273),
            .lcout(),
            .ltout(\Game_Inst.r_SM_Main_ns_i_i_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_1_LC_6_12_3 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_1_LC_6_12_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_SM_Main_1_LC_6_12_3 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \Game_Inst.r_SM_Main_1_LC_6_12_3  (
            .in0(N__7397),
            .in1(N__7680),
            .in2(N__4607),
            .in3(N__5264),
            .lcout(\Game_Inst.r_SM_MainZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8243),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_DV_RNIP6I59_LC_6_12_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_DV_RNIP6I59_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Button_DV_RNIP6I59_LC_6_12_6 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \Game_Inst.r_Button_DV_RNIP6I59_LC_6_12_6  (
            .in0(N__4598),
            .in1(N__5375),
            .in2(_gnd_net_),
            .in3(N__4580),
            .lcout(\Game_Inst.N_260_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_RNIJ6T62_12_LC_7_3_3 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_RNIJ6T62_12_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_Count_RNIJ6T62_12_LC_7_3_3 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \Debounce_SW4.r_Count_RNIJ6T62_12_LC_7_3_3  (
            .in0(N__5029),
            .in1(N__4760),
            .in2(N__5006),
            .in3(N__4766),
            .lcout(),
            .ltout(\Debounce_SW4.N_181_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_State_e_0_RNISK6T2_LC_7_3_4 .C_ON=1'b0;
    defparam \Debounce_SW4.r_State_e_0_RNISK6T2_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_State_e_0_RNISK6T2_LC_7_3_4 .LUT_INIT=16'b1111100110011001;
    LogicCell40 \Debounce_SW4.r_State_e_0_RNISK6T2_LC_7_3_4  (
            .in0(N__5438),
            .in1(N__8313),
            .in2(N__4781),
            .in3(N__5474),
            .lcout(\Debounce_SW4.N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_RNI55EK_4_LC_7_4_2 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_RNI55EK_4_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_Count_RNI55EK_4_LC_7_4_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Debounce_SW4.r_Count_RNI55EK_4_LC_7_4_2  (
            .in0(N__4846),
            .in1(N__4861),
            .in2(_gnd_net_),
            .in3(N__4876),
            .lcout(\Debounce_SW4.N_149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_RNIEO7R_1_LC_7_4_3 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_RNIEO7R_1_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_Count_RNIEO7R_1_LC_7_4_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW4.r_Count_RNIEO7R_1_LC_7_4_3  (
            .in0(N__4909),
            .in1(N__4730),
            .in2(N__4895),
            .in3(N__4707),
            .lcout(\Debounce_SW4.un9_r_count_10 ),
            .ltout(\Debounce_SW4.un9_r_count_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_RNIC1GM1_7_LC_7_4_4 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_RNIC1GM1_7_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_Count_RNIC1GM1_7_LC_7_4_4 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \Debounce_SW4.r_Count_RNIC1GM1_7_LC_7_4_4  (
            .in0(_gnd_net_),
            .in1(N__4830),
            .in2(N__4769),
            .in3(N__4750),
            .lcout(\Debounce_SW4.N_288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_RNISL0F_10_LC_7_4_5 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_RNISL0F_10_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_Count_RNISL0F_10_LC_7_4_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Debounce_SW4.r_Count_RNISL0F_10_LC_7_4_5  (
            .in0(N__5069),
            .in1(N__4799),
            .in2(N__5051),
            .in3(N__4813),
            .lcout(\Debounce_SW4.N_158 ),
            .ltout(\Debounce_SW4.N_158_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_State_e_0_RNO_0_LC_7_4_6 .C_ON=1'b0;
    defparam \Debounce_SW4.r_State_e_0_RNO_0_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_State_e_0_RNO_0_LC_7_4_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Debounce_SW4.r_State_e_0_RNO_0_LC_7_4_6  (
            .in0(N__5030),
            .in1(N__5005),
            .in2(N__4754),
            .in3(N__4831),
            .lcout(),
            .ltout(\Debounce_SW4.un9_r_count_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_State_e_0_RNO_LC_7_4_7 .C_ON=1'b0;
    defparam \Debounce_SW4.r_State_e_0_RNO_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_State_e_0_RNO_LC_7_4_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Debounce_SW4.r_State_e_0_RNO_LC_7_4_7  (
            .in0(N__4751),
            .in1(N__4742),
            .in2(N__4736),
            .in3(N__5473),
            .lcout(\Debounce_SW4.r_State_e_0_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.un2_r_count_cry_1_c_LC_7_5_0 .C_ON=1'b1;
    defparam \Debounce_SW4.un2_r_count_cry_1_c_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.un2_r_count_cry_1_c_LC_7_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Debounce_SW4.un2_r_count_cry_1_c_LC_7_5_0  (
            .in0(_gnd_net_),
            .in1(N__4731),
            .in2(N__4712),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_5_0_),
            .carryout(\Debounce_SW4.un2_r_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_2_LC_7_5_1 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_2_LC_7_5_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_2_LC_7_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_2_LC_7_5_1  (
            .in0(_gnd_net_),
            .in1(N__4910),
            .in2(_gnd_net_),
            .in3(N__4898),
            .lcout(\Debounce_SW4.r_CountZ0Z_2 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_1 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_2 ),
            .clk(N__8246),
            .ce(),
            .sr(N__4964));
    defparam \Debounce_SW4.r_Count_3_LC_7_5_2 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_3_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_3_LC_7_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_3_LC_7_5_2  (
            .in0(_gnd_net_),
            .in1(N__4894),
            .in2(_gnd_net_),
            .in3(N__4880),
            .lcout(\Debounce_SW4.r_CountZ0Z_3 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_2 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_3 ),
            .clk(N__8246),
            .ce(),
            .sr(N__4964));
    defparam \Debounce_SW4.r_Count_4_LC_7_5_3 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_4_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_4_LC_7_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_4_LC_7_5_3  (
            .in0(_gnd_net_),
            .in1(N__4877),
            .in2(_gnd_net_),
            .in3(N__4865),
            .lcout(\Debounce_SW4.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_3 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_4 ),
            .clk(N__8246),
            .ce(),
            .sr(N__4964));
    defparam \Debounce_SW4.r_Count_5_LC_7_5_4 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_5_LC_7_5_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_5_LC_7_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_5_LC_7_5_4  (
            .in0(_gnd_net_),
            .in1(N__4862),
            .in2(_gnd_net_),
            .in3(N__4850),
            .lcout(\Debounce_SW4.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_4 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_5 ),
            .clk(N__8246),
            .ce(),
            .sr(N__4964));
    defparam \Debounce_SW4.r_Count_6_LC_7_5_5 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_6_LC_7_5_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_6_LC_7_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_6_LC_7_5_5  (
            .in0(_gnd_net_),
            .in1(N__4847),
            .in2(_gnd_net_),
            .in3(N__4835),
            .lcout(\Debounce_SW4.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_5 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_6 ),
            .clk(N__8246),
            .ce(),
            .sr(N__4964));
    defparam \Debounce_SW4.r_Count_7_LC_7_5_6 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_7_LC_7_5_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_7_LC_7_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_7_LC_7_5_6  (
            .in0(_gnd_net_),
            .in1(N__4832),
            .in2(_gnd_net_),
            .in3(N__4817),
            .lcout(\Debounce_SW4.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_6 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_7 ),
            .clk(N__8246),
            .ce(),
            .sr(N__4964));
    defparam \Debounce_SW4.r_Count_8_LC_7_5_7 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_8_LC_7_5_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_8_LC_7_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_8_LC_7_5_7  (
            .in0(_gnd_net_),
            .in1(N__4814),
            .in2(_gnd_net_),
            .in3(N__4802),
            .lcout(\Debounce_SW4.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_7 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_8 ),
            .clk(N__8246),
            .ce(),
            .sr(N__4964));
    defparam \Debounce_SW4.r_Count_9_LC_7_6_0 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_9_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_9_LC_7_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_9_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__4798),
            .in2(_gnd_net_),
            .in3(N__4784),
            .lcout(\Debounce_SW4.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_7_6_0_),
            .carryout(\Debounce_SW4.un2_r_count_cry_9 ),
            .clk(N__8239),
            .ce(),
            .sr(N__4966));
    defparam \Debounce_SW4.r_Count_10_LC_7_6_1 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_10_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_10_LC_7_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_10_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__5068),
            .in2(_gnd_net_),
            .in3(N__5054),
            .lcout(\Debounce_SW4.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_9 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_10 ),
            .clk(N__8239),
            .ce(),
            .sr(N__4966));
    defparam \Debounce_SW4.r_Count_11_LC_7_6_2 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_11_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_11_LC_7_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_11_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__5047),
            .in2(_gnd_net_),
            .in3(N__5033),
            .lcout(\Debounce_SW4.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_10 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_11 ),
            .clk(N__8239),
            .ce(),
            .sr(N__4966));
    defparam \Debounce_SW4.r_Count_12_LC_7_6_3 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_12_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_12_LC_7_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_12_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__5028),
            .in2(_gnd_net_),
            .in3(N__5009),
            .lcout(\Debounce_SW4.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_11 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_12 ),
            .clk(N__8239),
            .ce(),
            .sr(N__4966));
    defparam \Debounce_SW4.r_Count_13_LC_7_6_4 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_13_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_13_LC_7_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_13_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(N__5001),
            .in2(_gnd_net_),
            .in3(N__4982),
            .lcout(\Debounce_SW4.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_12 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_13 ),
            .clk(N__8239),
            .ce(),
            .sr(N__4966));
    defparam \Debounce_SW4.r_Count_14_LC_7_6_5 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_14_LC_7_6_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_14_LC_7_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_14_LC_7_6_5  (
            .in0(_gnd_net_),
            .in1(N__5500),
            .in2(_gnd_net_),
            .in3(N__4979),
            .lcout(\Debounce_SW4.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_13 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_14 ),
            .clk(N__8239),
            .ce(),
            .sr(N__4966));
    defparam \Debounce_SW4.r_Count_15_LC_7_6_6 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_15_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_15_LC_7_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_15_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(N__5534),
            .in2(_gnd_net_),
            .in3(N__4976),
            .lcout(\Debounce_SW4.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_14 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_15 ),
            .clk(N__8239),
            .ce(),
            .sr(N__4966));
    defparam \Debounce_SW4.r_Count_16_LC_7_6_7 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_16_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_16_LC_7_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_16_LC_7_6_7  (
            .in0(_gnd_net_),
            .in1(N__5521),
            .in2(_gnd_net_),
            .in3(N__4973),
            .lcout(\Debounce_SW4.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Debounce_SW4.un2_r_count_cry_15 ),
            .carryout(\Debounce_SW4.un2_r_count_cry_16 ),
            .clk(N__8239),
            .ce(),
            .sr(N__4966));
    defparam \Debounce_SW4.r_Count_17_LC_7_7_0 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_17_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_17_LC_7_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Debounce_SW4.r_Count_17_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__5486),
            .in2(_gnd_net_),
            .in3(N__4970),
            .lcout(\Debounce_SW4.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8234),
            .ce(),
            .sr(N__4967));
    defparam \Debounce_SW1.r_Count_RNI2KFA_1_LC_7_8_1 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_RNI2KFA_1_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_RNI2KFA_1_LC_7_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW1.r_Count_RNI2KFA_1_LC_7_8_1  (
            .in0(N__4949),
            .in1(N__5895),
            .in2(N__4931),
            .in3(N__5873),
            .lcout(\Debounce_SW1.un9_r_count_10 ),
            .ltout(\Debounce_SW1.un9_r_count_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_RNIKOVK_7_LC_7_8_2 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_RNIKOVK_7_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_RNIKOVK_7_LC_7_8_2 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \Debounce_SW1.r_Count_RNIKOVK_7_LC_7_8_2  (
            .in0(_gnd_net_),
            .in1(N__5761),
            .in2(N__5126),
            .in3(N__5836),
            .lcout(),
            .ltout(\Debounce_SW1.N_285_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_RNI9B4K1_12_LC_7_8_3 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_RNI9B4K1_12_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_RNI9B4K1_12_LC_7_8_3 .LUT_INIT=16'b1110111011101010;
    LogicCell40 \Debounce_SW1.r_Count_RNI9B4K1_12_LC_7_8_3  (
            .in0(N__5782),
            .in1(N__5812),
            .in2(N__5123),
            .in3(N__5710),
            .lcout(),
            .ltout(\Debounce_SW1.N_184_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_State_e_0_RNI0MBO2_LC_7_8_4 .C_ON=1'b0;
    defparam \Debounce_SW1.r_State_e_0_RNI0MBO2_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_State_e_0_RNI0MBO2_LC_7_8_4 .LUT_INIT=16'b1110110010110011;
    LogicCell40 \Debounce_SW1.r_State_e_0_RNI0MBO2_LC_7_8_4  (
            .in0(N__5728),
            .in1(N__6758),
            .in2(N__5120),
            .in3(N__7105),
            .lcout(\Debounce_SW1.N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_4_RNIG59R_LC_7_8_7 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_4_RNIG59R_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Switch_4_RNIG59R_LC_7_8_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \Game_Inst.r_Switch_4_RNIG59R_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(N__5696),
            .in2(_gnd_net_),
            .in3(N__8331),
            .lcout(\Game_Inst.N_167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Toggle_LC_7_9_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Toggle_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Toggle_LC_7_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Toggle_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5647),
            .lcout(\Game_Inst.r_ToggleZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8235),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_ID_0_LC_7_9_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_ID_0_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Button_ID_0_LC_7_9_3 .LUT_INIT=16'b0000000011110100;
    LogicCell40 \Game_Inst.r_Button_ID_0_LC_7_9_3  (
            .in0(N__5098),
            .in1(N__8287),
            .in2(N__5087),
            .in3(N__5683),
            .lcout(\Game_Inst.r_Button_IDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8235),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_2_RNICD4F_LC_7_9_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_2_RNICD4F_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Switch_2_RNICD4F_LC_7_9_4 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \Game_Inst.r_Switch_2_RNICD4F_LC_7_9_4  (
            .in0(N__8051),
            .in1(N__5690),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Game_Inst.N_255 ),
            .ltout(\Game_Inst.N_255_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_DV_LC_7_9_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_DV_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Button_DV_LC_7_9_5 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \Game_Inst.r_Button_DV_LC_7_9_5  (
            .in0(N__5097),
            .in1(N__8286),
            .in2(N__5102),
            .in3(N__5682),
            .lcout(\Game_Inst.r_Button_DVZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8235),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_ID_1_LC_7_9_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_ID_1_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Button_ID_1_LC_7_9_6 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \Game_Inst.r_Button_ID_1_LC_7_9_6  (
            .in0(N__5684),
            .in1(N__5099),
            .in2(N__8291),
            .in3(N__5086),
            .lcout(\Game_Inst.r_Button_IDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8235),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_0_RNIFS911_1_LC_7_10_0 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_0_RNIFS911_1_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_0_RNIFS911_1_LC_7_10_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Game_Inst.r_Pattern_0_RNIFS911_1_LC_7_10_0  (
            .in0(N__5936),
            .in1(N__5336),
            .in2(_gnd_net_),
            .in3(N__5927),
            .lcout(),
            .ltout(\Game_Inst.r_Pattern_0_RNIFS911Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNIHD922_1_LC_7_10_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNIHD922_1_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNIHD922_1_LC_7_10_1 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \Game_Inst.r_Index_RNIHD922_1_LC_7_10_1  (
            .in0(N__5211),
            .in1(N__5244),
            .in2(N__5219),
            .in3(N__5180),
            .lcout(),
            .ltout(\Game_Inst.un6_r_button_dv_7_i_m2_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNIRNF03_2_LC_7_10_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNIRNF03_2_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNIRNF03_2_LC_7_10_2 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \Game_Inst.r_Index_RNIRNF03_2_LC_7_10_2  (
            .in0(N__5144),
            .in1(N__5212),
            .in2(N__5189),
            .in3(N__5138),
            .lcout(\Game_Inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_3_RNIH6ML_0_LC_7_10_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_3_RNIH6ML_0_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_3_RNIH6ML_0_LC_7_10_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Game_Inst.r_Pattern_3_RNIH6ML_0_LC_7_10_3  (
            .in0(N__5334),
            .in1(N__5915),
            .in2(_gnd_net_),
            .in3(N__5909),
            .lcout(\Game_Inst.r_Pattern_3_RNIH6MLZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_3_RNIJ8ML_1_LC_7_10_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_3_RNIJ8ML_1_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_3_RNIJ8ML_1_LC_7_10_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Game_Inst.r_Pattern_3_RNIJ8ML_1_LC_7_10_4  (
            .in0(N__5966),
            .in1(N__5333),
            .in2(_gnd_net_),
            .in3(N__5972),
            .lcout(\Game_Inst.r_Pattern_3_RNIJ8MLZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_0_0_LC_7_10_5 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_0_0_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_0_0_LC_7_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_0_0_LC_7_10_5  (
            .in0(N__5984),
            .in1(N__5132),
            .in2(N__5174),
            .in3(N__7299),
            .lcout(\Game_Inst.r_SM_Main_ns_i_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_6_RNIR0FE_1_LC_7_10_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_6_RNIR0FE_1_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_6_RNIR0FE_1_LC_7_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Game_Inst.r_Pattern_6_RNIR0FE_1_LC_7_10_6  (
            .in0(N__5337),
            .in1(N__5921),
            .in2(_gnd_net_),
            .in3(N__6086),
            .lcout(\Game_Inst.r_Pattern_6_RNIR0FEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_4_RNINK2A_1_LC_7_10_7 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_4_RNINK2A_1_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_4_RNINK2A_1_LC_7_10_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Game_Inst.r_Pattern_4_RNINK2A_1_LC_7_10_7  (
            .in0(N__5335),
            .in1(N__6080),
            .in2(_gnd_net_),
            .in3(N__6116),
            .lcout(\Game_Inst.r_Pattern_4_RNINK2AZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_3_0_LC_7_11_0 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_3_0_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_3_0_LC_7_11_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_3_0_LC_7_11_0  (
            .in0(N__6042),
            .in1(N__7467),
            .in2(N__7576),
            .in3(N__7387),
            .lcout(\Game_Inst.N_266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI9A2A_0_0_LC_7_11_1 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI9A2A_0_0_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI9A2A_0_0_LC_7_11_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Game_Inst.r_SM_Main_RNI9A2A_0_0_LC_7_11_1  (
            .in0(N__7386),
            .in1(N__7540),
            .in2(_gnd_net_),
            .in3(N__7686),
            .lcout(\Game_Inst.r_SM_Main_d_6 ),
            .ltout(\Game_Inst.r_SM_Main_d_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_DV_RNIP62M_LC_7_11_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_DV_RNIP62M_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Button_DV_RNIP62M_LC_7_11_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Game_Inst.r_Button_DV_RNIP62M_LC_7_11_2  (
            .in0(N__5371),
            .in1(N__8047),
            .in2(N__5348),
            .in3(N__7113),
            .lcout(\Game_Inst.r_Score_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_4_RNILI2A_0_LC_7_11_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_4_RNILI2A_0_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_4_RNILI2A_0_LC_7_11_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Game_Inst.r_Pattern_4_RNILI2A_0_LC_7_11_3  (
            .in0(N__5978),
            .in1(N__6110),
            .in2(_gnd_net_),
            .in3(N__5330),
            .lcout(\Game_Inst.r_Pattern_4_RNILI2AZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_2_LC_7_11_4 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_2_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_2_LC_7_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_2_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5959),
            .lcout(\Game_Inst.w_LFSR_Data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8245),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_3_1_LC_7_12_0 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_3_1_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_3_1_LC_7_12_0 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_3_1_LC_7_12_0  (
            .in0(N__6043),
            .in1(N__7393),
            .in2(N__7593),
            .in3(N__7696),
            .lcout(\Game_Inst.N_259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_0_2_LC_7_12_5 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_0_2_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_0_2_LC_7_12_5 .LUT_INIT=16'b0000010001011111;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_0_2_LC_7_12_5  (
            .in0(N__7697),
            .in1(N__6044),
            .in2(N__7415),
            .in3(N__7566),
            .lcout(),
            .ltout(\Game_Inst.r_SM_Main_ns_i_0_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_2_LC_7_12_6 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_2_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_SM_Main_2_LC_7_12_6 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \Game_Inst.r_SM_Main_2_LC_7_12_6  (
            .in0(N__7567),
            .in1(N__7483),
            .in2(N__5267),
            .in3(N__5263),
            .lcout(\Game_Inst.r_SM_MainZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8249),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.un2_r_count_cry_1_c_LC_7_13_0 .C_ON=1'b1;
    defparam \Debounce_SW2.un2_r_count_cry_1_c_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.un2_r_count_cry_1_c_LC_7_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Debounce_SW2.un2_r_count_cry_1_c_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__6437),
            .in2(N__6461),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\Debounce_SW2.un2_r_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_2_LC_7_13_1 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_2_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_2_LC_7_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_2_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__6557),
            .in2(_gnd_net_),
            .in3(N__5252),
            .lcout(\Debounce_SW2.r_CountZ0Z_2 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_1 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_2 ),
            .clk(N__8256),
            .ce(),
            .sr(N__6413));
    defparam \Debounce_SW2.r_Count_3_LC_7_13_2 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_3_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_3_LC_7_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_3_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__6544),
            .in2(_gnd_net_),
            .in3(N__5402),
            .lcout(\Debounce_SW2.r_CountZ0Z_3 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_2 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_3 ),
            .clk(N__8256),
            .ce(),
            .sr(N__6413));
    defparam \Debounce_SW2.r_Count_4_LC_7_13_3 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_4_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_4_LC_7_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_4_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__6137),
            .in2(_gnd_net_),
            .in3(N__5399),
            .lcout(\Debounce_SW2.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_3 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_4 ),
            .clk(N__8256),
            .ce(),
            .sr(N__6413));
    defparam \Debounce_SW2.r_Count_5_LC_7_13_4 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_5_LC_7_13_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_5_LC_7_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_5_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__6149),
            .in2(_gnd_net_),
            .in3(N__5396),
            .lcout(\Debounce_SW2.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_4 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_5 ),
            .clk(N__8256),
            .ce(),
            .sr(N__6413));
    defparam \Debounce_SW2.r_Count_6_LC_7_13_5 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_6_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_6_LC_7_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_6_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__6161),
            .in2(_gnd_net_),
            .in3(N__5393),
            .lcout(\Debounce_SW2.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_5 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_6 ),
            .clk(N__8256),
            .ce(),
            .sr(N__6413));
    defparam \Debounce_SW2.r_Count_7_LC_7_13_6 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_7_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_7_LC_7_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_7_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__6581),
            .in2(_gnd_net_),
            .in3(N__5390),
            .lcout(\Debounce_SW2.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_6 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_7 ),
            .clk(N__8256),
            .ce(),
            .sr(N__6413));
    defparam \Debounce_SW2.r_Count_8_LC_7_13_7 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_8_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_8_LC_7_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_8_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__6221),
            .in2(_gnd_net_),
            .in3(N__5387),
            .lcout(\Debounce_SW2.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_7 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_8 ),
            .clk(N__8256),
            .ce(),
            .sr(N__6413));
    defparam \Debounce_SW2.r_Count_9_LC_7_14_0 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_9_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_9_LC_7_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_9_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__6248),
            .in2(_gnd_net_),
            .in3(N__5384),
            .lcout(\Debounce_SW2.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\Debounce_SW2.un2_r_count_cry_9 ),
            .clk(N__8262),
            .ce(),
            .sr(N__6411));
    defparam \Debounce_SW2.r_Count_10_LC_7_14_1 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_10_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_10_LC_7_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_10_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__6260),
            .in2(_gnd_net_),
            .in3(N__5381),
            .lcout(\Debounce_SW2.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_9 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_10 ),
            .clk(N__8262),
            .ce(),
            .sr(N__6411));
    defparam \Debounce_SW2.r_Count_11_LC_7_14_2 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_11_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_11_LC_7_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_11_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__6235),
            .in2(_gnd_net_),
            .in3(N__5378),
            .lcout(\Debounce_SW2.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_10 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_11 ),
            .clk(N__8262),
            .ce(),
            .sr(N__6411));
    defparam \Debounce_SW2.r_Count_12_LC_7_14_3 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_12_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_12_LC_7_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_12_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__6188),
            .in2(_gnd_net_),
            .in3(N__5456),
            .lcout(\Debounce_SW2.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_11 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_12 ),
            .clk(N__8262),
            .ce(),
            .sr(N__6411));
    defparam \Debounce_SW2.r_Count_13_LC_7_14_4 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_13_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_13_LC_7_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_13_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__6208),
            .in2(_gnd_net_),
            .in3(N__5453),
            .lcout(\Debounce_SW2.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_12 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_13 ),
            .clk(N__8262),
            .ce(),
            .sr(N__6411));
    defparam \Debounce_SW2.r_Count_14_LC_7_14_5 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_14_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_14_LC_7_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_14_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__6482),
            .in2(_gnd_net_),
            .in3(N__5450),
            .lcout(\Debounce_SW2.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_13 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_14 ),
            .clk(N__8262),
            .ce(),
            .sr(N__6411));
    defparam \Debounce_SW2.r_Count_15_LC_7_14_6 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_15_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_15_LC_7_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_15_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__6509),
            .in2(_gnd_net_),
            .in3(N__5447),
            .lcout(\Debounce_SW2.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_14 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_15 ),
            .clk(N__8262),
            .ce(),
            .sr(N__6411));
    defparam \Debounce_SW2.r_Count_16_LC_7_14_7 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_16_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_16_LC_7_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_16_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(N__6521),
            .in2(_gnd_net_),
            .in3(N__5444),
            .lcout(\Debounce_SW2.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Debounce_SW2.un2_r_count_cry_15 ),
            .carryout(\Debounce_SW2.un2_r_count_cry_16 ),
            .clk(N__8262),
            .ce(),
            .sr(N__6411));
    defparam \Debounce_SW2.r_Count_17_LC_7_15_0 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_17_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_17_LC_7_15_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Debounce_SW2.r_Count_17_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__6496),
            .in2(_gnd_net_),
            .in3(N__5441),
            .lcout(\Debounce_SW2.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8265),
            .ce(),
            .sr(N__6410));
    defparam \Debounce_SW4.r_State_e_0_LC_8_3_0 .C_ON=1'b0;
    defparam \Debounce_SW4.r_State_e_0_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_State_e_0_LC_8_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Debounce_SW4.r_State_e_0_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5434),
            .lcout(w_Switch_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8263),
            .ce(N__5411),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_1_LC_8_4_2 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_1_LC_8_4_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_1_LC_8_4_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Debounce_SW3.r_Count_1_LC_8_4_2  (
            .in0(N__6395),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6373),
            .lcout(\Debounce_SW3.r_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8258),
            .ce(),
            .sr(N__6776));
    defparam \Debounce_SW3.r_Count_0_LC_8_4_5 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_0_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_0_LC_8_4_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Debounce_SW3.r_Count_0_LC_8_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6394),
            .lcout(\Debounce_SW3.r_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8258),
            .ce(),
            .sr(N__6776));
    defparam \Debounce_SW3.r_Count_RNIACA_1_LC_8_5_3 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_RNIACA_1_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_RNIACA_1_LC_8_5_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW3.r_Count_RNIACA_1_LC_8_5_3  (
            .in0(N__6352),
            .in1(N__6369),
            .in2(N__6338),
            .in3(N__6392),
            .lcout(\Debounce_SW3.un9_r_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_RNI248_4_LC_8_5_5 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_RNI248_4_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_RNI248_4_LC_8_5_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Debounce_SW3.r_Count_RNI248_4_LC_8_5_5  (
            .in0(N__6697),
            .in1(N__6712),
            .in2(_gnd_net_),
            .in3(N__6727),
            .lcout(\Debounce_SW3.N_148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_RNI58AB_12_LC_8_6_0 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_RNI58AB_12_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_RNI58AB_12_LC_8_6_0 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \Debounce_SW3.r_Count_RNI58AB_12_LC_8_6_0  (
            .in0(N__6597),
            .in1(N__5576),
            .in2(N__6866),
            .in3(N__5567),
            .lcout(\Debounce_SW3.N_182 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_RNIO7D5_8_LC_8_6_1 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_RNIO7D5_8_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_RNIO7D5_8_LC_8_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Debounce_SW3.r_Count_RNIO7D5_8_LC_8_6_1  (
            .in0(N__6635),
            .in1(N__6649),
            .in2(N__6617),
            .in3(N__6664),
            .lcout(\Debounce_SW3.N_159 ),
            .ltout(\Debounce_SW3.N_159_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_State_e_0_RNO_0_LC_8_6_2 .C_ON=1'b0;
    defparam \Debounce_SW3.r_State_e_0_RNO_0_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_State_e_0_RNO_0_LC_8_6_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Debounce_SW3.r_State_e_0_RNO_0_LC_8_6_2  (
            .in0(N__6598),
            .in1(N__6864),
            .in2(N__5570),
            .in3(N__6682),
            .lcout(\Debounce_SW3.un9_r_count_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_RNI49L_7_LC_8_6_3 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_RNI49L_7_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_RNI49L_7_LC_8_6_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \Debounce_SW3.r_Count_RNI49L_7_LC_8_6_3  (
            .in0(N__6681),
            .in1(N__5554),
            .in2(_gnd_net_),
            .in3(N__5542),
            .lcout(\Debounce_SW3.N_287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_RNIUQFA_17_LC_8_6_4 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_RNIUQFA_17_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_RNIUQFA_17_LC_8_6_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW3.r_Count_RNIUQFA_17_LC_8_6_4  (
            .in0(N__6811),
            .in1(N__6826),
            .in2(N__6794),
            .in3(N__6841),
            .lcout(\Debounce_SW3.r_count15_i_a2_0 ),
            .ltout(\Debounce_SW3.r_count15_i_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_State_e_0_RNO_LC_8_6_5 .C_ON=1'b0;
    defparam \Debounce_SW3.r_State_e_0_RNO_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_State_e_0_RNO_LC_8_6_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Debounce_SW3.r_State_e_0_RNO_LC_8_6_5  (
            .in0(N__5561),
            .in1(N__5555),
            .in2(N__5546),
            .in3(N__5543),
            .lcout(\Debounce_SW3.r_State_e_0_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_RNI2BP2_17_LC_8_6_6 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_RNI2BP2_17_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_Count_RNI2BP2_17_LC_8_6_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW4.r_Count_RNI2BP2_17_LC_8_6_6  (
            .in0(N__5533),
            .in1(N__5522),
            .in2(N__5507),
            .in3(N__5485),
            .lcout(\Debounce_SW4.r_count15_i_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_1_LC_8_7_4 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_1_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_1_LC_8_7_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Debounce_SW1.r_Count_1_LC_8_7_4  (
            .in0(N__5878),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5899),
            .lcout(\Debounce_SW1.r_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8240),
            .ce(),
            .sr(N__5855));
    defparam \Debounce_SW1.r_Count_0_LC_8_7_7 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_0_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_0_LC_8_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Debounce_SW1.r_Count_0_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5877),
            .lcout(\Debounce_SW1.r_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8240),
            .ce(),
            .sr(N__5855));
    defparam \Debounce_SW1.r_State_e_0_RNO_0_LC_8_8_0 .C_ON=1'b0;
    defparam \Debounce_SW1.r_State_e_0_RNO_0_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_State_e_0_RNO_0_LC_8_8_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Debounce_SW1.r_State_e_0_RNO_0_LC_8_8_0  (
            .in0(N__5837),
            .in1(N__5813),
            .in2(N__5789),
            .in3(N__5762),
            .lcout(),
            .ltout(\Debounce_SW1.un9_r_count_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_State_e_0_RNO_LC_8_8_1 .C_ON=1'b0;
    defparam \Debounce_SW1.r_State_e_0_RNO_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_State_e_0_RNO_LC_8_8_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Debounce_SW1.r_State_e_0_RNO_LC_8_8_1  (
            .in0(N__5738),
            .in1(N__5732),
            .in2(N__5714),
            .in3(N__5711),
            .lcout(\Debounce_SW1.r_State_e_0_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_4_LC_8_8_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_4_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Switch_4_LC_8_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Switch_4_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8332),
            .lcout(\Game_Inst.r_SwitchZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8229),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_2_LC_8_9_0 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_2_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Switch_2_LC_8_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Switch_2_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8052),
            .lcout(\Game_Inst.r_SwitchZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8241),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_1_RNIA12H_LC_8_9_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_1_RNIA12H_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Switch_1_RNIA12H_LC_8_9_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Game_Inst.r_Switch_1_RNIA12H_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__5672),
            .in2(_gnd_net_),
            .in3(N__7093),
            .lcout(\Game_Inst.r_Switch_1_RNIA12HZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_1_LC_8_9_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_1_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Switch_1_LC_8_9_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Game_Inst.r_Switch_1_LC_8_9_2  (
            .in0(N__7094),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Game_Inst.r_SwitchZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8241),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_4_0_LC_8_9_3 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_4_0_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_4_0_LC_8_9_3 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_4_0_LC_8_9_3  (
            .in0(N__5657),
            .in1(N__5592),
            .in2(_gnd_net_),
            .in3(N__7599),
            .lcout(),
            .ltout(\Game_Inst.N_208_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_2_0_LC_8_9_4 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_2_0_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_2_0_LC_8_9_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_2_0_LC_8_9_4  (
            .in0(N__7468),
            .in1(N__7417),
            .in2(N__5987),
            .in3(N__7698),
            .lcout(\Game_Inst.N_264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_5_0_LC_8_10_0 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_5_0_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_5_0_LC_8_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_5_0_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6992),
            .lcout(\Game_Inst.r_Pattern_5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8247),
            .ce(N__6074),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_3_1_LC_8_10_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_3_1_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_3_1_LC_8_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_3_1_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6029),
            .lcout(\Game_Inst.r_Pattern_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8247),
            .ce(N__6074),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_2_1_LC_8_10_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_2_1_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_2_1_LC_8_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_2_1_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6320),
            .lcout(\Game_Inst.r_Pattern_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8247),
            .ce(N__6074),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_0_1_LC_8_10_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_0_1_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_0_1_LC_8_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_0_1_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5960),
            .lcout(\Game_Inst.r_Pattern_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8247),
            .ce(N__6074),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_1_1_LC_8_10_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_1_1_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_1_1_LC_8_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_1_1_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6305),
            .lcout(\Game_Inst.r_Pattern_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8247),
            .ce(N__6074),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_6_1_LC_8_10_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_6_1_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_6_1_LC_8_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_6_1_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7003),
            .lcout(\Game_Inst.r_Pattern_6Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8247),
            .ce(N__6074),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_2_0_LC_8_10_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_2_0_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_2_0_LC_8_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_2_0_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6290),
            .lcout(\Game_Inst.r_Pattern_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8247),
            .ce(N__6074),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_3_0_LC_8_11_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_3_0_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_3_0_LC_8_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_3_0_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5999),
            .lcout(\Game_Inst.r_Pattern_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8250),
            .ce(N__6066),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_4_1_LC_8_11_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_4_1_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_4_1_LC_8_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_4_1_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7174),
            .lcout(\Game_Inst.r_Pattern_4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8250),
            .ce(N__6066),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_4_0_LC_8_11_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_4_0_LC_8_11_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_4_0_LC_8_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_4_0_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7187),
            .lcout(\Game_Inst.r_Pattern_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8250),
            .ce(N__6066),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_7_1_LC_8_11_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_7_1_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_7_1_LC_8_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_7_1_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6104),
            .lcout(\Game_Inst.r_Pattern_7Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8250),
            .ce(N__6066),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_5_1_LC_8_11_7 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_5_1_LC_8_11_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_5_1_LC_8_11_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \Game_Inst.r_Pattern_5_1_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__7040),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Game_Inst.r_Pattern_5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8250),
            .ce(N__6066),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_17_6_0__m5_0_o2_LC_8_12_0 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_17_6_0__m5_0_o2_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \Scoreboard.r_Hex_Encoding_17_6_0__m5_0_o2_LC_8_12_0 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \Scoreboard.r_Hex_Encoding_17_6_0__m5_0_o2_LC_8_12_0  (
            .in0(N__7210),
            .in1(N__7792),
            .in2(N__6913),
            .in3(N__7723),
            .lcout(N_143),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_7_LC_8_12_1 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_7_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_7_LC_8_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_7_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5998),
            .lcout(\Game_Inst.w_LFSR_Data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8257),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_8_LC_8_12_2 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_8_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_8_LC_8_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_8_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6025),
            .lcout(\Game_Inst.w_LFSR_Data_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8257),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_3_LC_8_12_3 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_3_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_3_LC_8_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_3_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6013),
            .lcout(\Game_Inst.w_LFSR_Data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8257),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_6_LC_8_12_4 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_6_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_6_LC_8_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_6_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6316),
            .lcout(\Game_Inst.w_LFSR_Data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8257),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_5_LC_8_12_5 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_5_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_5_LC_8_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_5_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6286),
            .lcout(\Game_Inst.w_LFSR_Data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8257),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_4_LC_8_12_7 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_4_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_4_LC_8_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_4_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6301),
            .lcout(\Game_Inst.w_LFSR_Data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8257),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_RNIN9NF3_12_LC_8_13_0 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_RNIN9NF3_12_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_RNIN9NF3_12_LC_8_13_0 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \Debounce_SW2.r_Count_RNIN9NF3_12_LC_8_13_0  (
            .in0(N__6186),
            .in1(N__6169),
            .in2(N__6209),
            .in3(N__6563),
            .lcout(),
            .ltout(\Debounce_SW2.N_183_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_State_e_0_RNIKLK44_LC_8_13_1 .C_ON=1'b0;
    defparam \Debounce_SW2.r_State_e_0_RNIKLK44_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_State_e_0_RNIKLK44_LC_8_13_1 .LUT_INIT=16'b1110110010110011;
    LogicCell40 \Debounce_SW2.r_State_e_0_RNIKLK44_LC_8_13_1  (
            .in0(N__6469),
            .in1(N__7160),
            .in2(N__6275),
            .in3(N__8016),
            .lcout(\Debounce_SW2.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_RNIKPPR_10_LC_8_13_2 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_RNIKPPR_10_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_RNIKPPR_10_LC_8_13_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Debounce_SW2.r_Count_RNIKPPR_10_LC_8_13_2  (
            .in0(N__6259),
            .in1(N__6247),
            .in2(N__6236),
            .in3(N__6220),
            .lcout(\Debounce_SW2.N_160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_State_e_0_RNO_0_LC_8_13_3 .C_ON=1'b0;
    defparam \Debounce_SW2.r_State_e_0_RNO_0_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_State_e_0_RNO_0_LC_8_13_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Debounce_SW2.r_State_e_0_RNO_0_LC_8_13_3  (
            .in0(N__6207),
            .in1(N__6187),
            .in2(N__6125),
            .in3(N__6580),
            .lcout(),
            .ltout(\Debounce_SW2.un9_r_count_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_State_e_0_RNO_LC_8_13_4 .C_ON=1'b0;
    defparam \Debounce_SW2.r_State_e_0_RNO_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_State_e_0_RNO_LC_8_13_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Debounce_SW2.r_State_e_0_RNO_LC_8_13_4  (
            .in0(N__6530),
            .in1(N__6470),
            .in2(N__6173),
            .in3(N__6170),
            .lcout(\Debounce_SW2.r_State_e_0_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_RNIV22S_4_LC_8_13_6 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_RNIV22S_4_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_RNIV22S_4_LC_8_13_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Debounce_SW2.r_Count_RNIV22S_4_LC_8_13_6  (
            .in0(N__6160),
            .in1(N__6148),
            .in2(_gnd_net_),
            .in3(N__6136),
            .lcout(\Debounce_SW2.N_147 ),
            .ltout(\Debounce_SW2.N_147_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_RNISGQA2_7_LC_8_13_7 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_RNISGQA2_7_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_RNISGQA2_7_LC_8_13_7 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \Debounce_SW2.r_Count_RNISGQA2_7_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__6579),
            .in2(N__6566),
            .in3(N__6529),
            .lcout(\Debounce_SW2.N_286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_RNI60D51_1_LC_8_14_2 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_RNI60D51_1_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_RNI60D51_1_LC_8_14_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW2.r_Count_RNI60D51_1_LC_8_14_2  (
            .in0(N__6556),
            .in1(N__6453),
            .in2(N__6545),
            .in3(N__6431),
            .lcout(\Debounce_SW2.un9_r_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_RNIQA6I_17_LC_8_14_6 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_RNIQA6I_17_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_RNIQA6I_17_LC_8_14_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW2.r_Count_RNIQA6I_17_LC_8_14_6  (
            .in0(N__6520),
            .in1(N__6508),
            .in2(N__6497),
            .in3(N__6481),
            .lcout(\Debounce_SW2.r_count15_i_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_1_LC_8_15_1 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_1_LC_8_15_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_1_LC_8_15_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Debounce_SW2.r_Count_1_LC_8_15_1  (
            .in0(N__6436),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6457),
            .lcout(\Debounce_SW2.r_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8267),
            .ce(),
            .sr(N__6412));
    defparam \Debounce_SW2.r_Count_0_LC_8_15_2 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_0_LC_8_15_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_0_LC_8_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Debounce_SW2.r_Count_0_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6435),
            .lcout(\Debounce_SW2.r_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8267),
            .ce(),
            .sr(N__6412));
    defparam \Debounce_SW3.un2_r_count_cry_1_c_LC_9_5_0 .C_ON=1'b1;
    defparam \Debounce_SW3.un2_r_count_cry_1_c_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.un2_r_count_cry_1_c_LC_9_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Debounce_SW3.un2_r_count_cry_1_c_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__6393),
            .in2(N__6374),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\Debounce_SW3.un2_r_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_2_LC_9_5_1 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_2_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_2_LC_9_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_2_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__6353),
            .in2(_gnd_net_),
            .in3(N__6341),
            .lcout(\Debounce_SW3.r_CountZ0Z_2 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_1 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_2 ),
            .clk(N__8260),
            .ce(),
            .sr(N__6775));
    defparam \Debounce_SW3.r_Count_3_LC_9_5_2 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_3_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_3_LC_9_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_3_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__6337),
            .in2(_gnd_net_),
            .in3(N__6323),
            .lcout(\Debounce_SW3.r_CountZ0Z_3 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_2 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_3 ),
            .clk(N__8260),
            .ce(),
            .sr(N__6775));
    defparam \Debounce_SW3.r_Count_4_LC_9_5_3 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_4_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_4_LC_9_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_4_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__6728),
            .in2(_gnd_net_),
            .in3(N__6716),
            .lcout(\Debounce_SW3.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_3 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_4 ),
            .clk(N__8260),
            .ce(),
            .sr(N__6775));
    defparam \Debounce_SW3.r_Count_5_LC_9_5_4 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_5_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_5_LC_9_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_5_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__6713),
            .in2(_gnd_net_),
            .in3(N__6701),
            .lcout(\Debounce_SW3.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_4 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_5 ),
            .clk(N__8260),
            .ce(),
            .sr(N__6775));
    defparam \Debounce_SW3.r_Count_6_LC_9_5_5 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_6_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_6_LC_9_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_6_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__6698),
            .in2(_gnd_net_),
            .in3(N__6686),
            .lcout(\Debounce_SW3.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_5 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_6 ),
            .clk(N__8260),
            .ce(),
            .sr(N__6775));
    defparam \Debounce_SW3.r_Count_7_LC_9_5_6 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_7_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_7_LC_9_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_7_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(N__6683),
            .in2(_gnd_net_),
            .in3(N__6668),
            .lcout(\Debounce_SW3.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_6 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_7 ),
            .clk(N__8260),
            .ce(),
            .sr(N__6775));
    defparam \Debounce_SW3.r_Count_8_LC_9_5_7 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_8_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_8_LC_9_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_8_LC_9_5_7  (
            .in0(_gnd_net_),
            .in1(N__6665),
            .in2(_gnd_net_),
            .in3(N__6653),
            .lcout(\Debounce_SW3.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_7 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_8 ),
            .clk(N__8260),
            .ce(),
            .sr(N__6775));
    defparam \Debounce_SW3.r_Count_9_LC_9_6_0 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_9_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_9_LC_9_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_9_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__6650),
            .in2(_gnd_net_),
            .in3(N__6638),
            .lcout(\Debounce_SW3.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\Debounce_SW3.un2_r_count_cry_9 ),
            .clk(N__8252),
            .ce(),
            .sr(N__6774));
    defparam \Debounce_SW3.r_Count_10_LC_9_6_1 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_10_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_10_LC_9_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_10_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__6634),
            .in2(_gnd_net_),
            .in3(N__6620),
            .lcout(\Debounce_SW3.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_9 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_10 ),
            .clk(N__8252),
            .ce(),
            .sr(N__6774));
    defparam \Debounce_SW3.r_Count_11_LC_9_6_2 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_11_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_11_LC_9_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_11_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__6616),
            .in2(_gnd_net_),
            .in3(N__6602),
            .lcout(\Debounce_SW3.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_10 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_11 ),
            .clk(N__8252),
            .ce(),
            .sr(N__6774));
    defparam \Debounce_SW3.r_Count_12_LC_9_6_3 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_12_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_12_LC_9_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_12_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(N__6599),
            .in2(_gnd_net_),
            .in3(N__6584),
            .lcout(\Debounce_SW3.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_11 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_12 ),
            .clk(N__8252),
            .ce(),
            .sr(N__6774));
    defparam \Debounce_SW3.r_Count_13_LC_9_6_4 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_13_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_13_LC_9_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_13_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__6865),
            .in2(_gnd_net_),
            .in3(N__6845),
            .lcout(\Debounce_SW3.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_12 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_13 ),
            .clk(N__8252),
            .ce(),
            .sr(N__6774));
    defparam \Debounce_SW3.r_Count_14_LC_9_6_5 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_14_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_14_LC_9_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_14_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(N__6842),
            .in2(_gnd_net_),
            .in3(N__6830),
            .lcout(\Debounce_SW3.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_13 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_14 ),
            .clk(N__8252),
            .ce(),
            .sr(N__6774));
    defparam \Debounce_SW3.r_Count_15_LC_9_6_6 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_15_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_15_LC_9_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_15_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__6827),
            .in2(_gnd_net_),
            .in3(N__6815),
            .lcout(\Debounce_SW3.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_14 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_15 ),
            .clk(N__8252),
            .ce(),
            .sr(N__6774));
    defparam \Debounce_SW3.r_Count_16_LC_9_6_7 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_16_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_16_LC_9_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_16_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(N__6812),
            .in2(_gnd_net_),
            .in3(N__6800),
            .lcout(\Debounce_SW3.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Debounce_SW3.un2_r_count_cry_15 ),
            .carryout(\Debounce_SW3.un2_r_count_cry_16 ),
            .clk(N__8252),
            .ce(),
            .sr(N__6774));
    defparam \Debounce_SW3.r_Count_17_LC_9_7_0 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_17_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_17_LC_9_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Debounce_SW3.r_Count_17_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__6790),
            .in2(_gnd_net_),
            .in3(N__6797),
            .lcout(\Debounce_SW3.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8248),
            .ce(),
            .sr(N__6773));
    defparam \Debounce_SW1.r_State_e_0_LC_9_8_5 .C_ON=1'b0;
    defparam \Debounce_SW1.r_State_e_0_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_State_e_0_LC_9_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Debounce_SW1.r_State_e_0_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6754),
            .lcout(w_Switch_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8236),
            .ce(N__6737),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI9A2A_0_LC_9_9_5 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI9A2A_0_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI9A2A_0_LC_9_9_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Game_Inst.r_SM_Main_RNI9A2A_0_LC_9_9_5  (
            .in0(N__7418),
            .in1(N__7600),
            .in2(_gnd_net_),
            .in3(N__7699),
            .lcout(\Game_Inst.N_338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_11_LC_9_10_0 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_11_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_11_LC_9_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_11_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6991),
            .lcout(\Game_Inst.w_LFSR_Data_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8251),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_12_LC_9_10_2 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_12_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_12_LC_9_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_12_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7039),
            .lcout(\Game_Inst.w_LFSR_Data_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8251),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_13_LC_9_10_4 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_13_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_13_LC_9_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_13_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7021),
            .lcout(\Game_Inst.w_LFSR_Data_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8251),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_10_LC_9_10_5 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_10_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_10_LC_9_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_10_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7175),
            .lcout(\Game_Inst.w_LFSR_Data_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8251),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Score_RNO_0_0_LC_9_11_0 .C_ON=1'b1;
    defparam \Game_Inst.r_Score_RNO_0_0_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Score_RNO_0_0_LC_9_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.r_Score_RNO_0_0_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__7730),
            .in2(N__6881),
            .in3(N__6880),
            .lcout(\Game_Inst.r_Score_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\Game_Inst.un1_r_Score_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.un1_r_Score_cry_0_THRU_LUT4_0_LC_9_11_1 .C_ON=1'b1;
    defparam \Game_Inst.un1_r_Score_cry_0_THRU_LUT4_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.un1_r_Score_cry_0_THRU_LUT4_0_LC_9_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.un1_r_Score_cry_0_THRU_LUT4_0_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__7801),
            .in2(_gnd_net_),
            .in3(N__6980),
            .lcout(\Game_Inst.un1_r_Score_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\Game_Inst.un1_r_Score_cry_0 ),
            .carryout(\Game_Inst.un1_r_Score_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Score_RNO_0_2_LC_9_11_2 .C_ON=1'b1;
    defparam \Game_Inst.r_Score_RNO_0_2_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Score_RNO_0_2_LC_9_11_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Game_Inst.r_Score_RNO_0_2_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7234),
            .in3(N__6977),
            .lcout(\Game_Inst.r_Score_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\Game_Inst.un1_r_Score_cry_1 ),
            .carryout(\Game_Inst.un1_r_Score_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Score_3_LC_9_11_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Score_3_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Score_3_LC_9_11_3 .LUT_INIT=16'b0010001100110010;
    LogicCell40 \Game_Inst.r_Score_3_LC_9_11_3  (
            .in0(N__7281),
            .in1(N__7315),
            .in2(N__6938),
            .in3(N__6974),
            .lcout(w_Score_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8259),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_0_sqmuxa_2_i_a2_2_LC_9_11_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_0_sqmuxa_2_i_a2_2_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_0_sqmuxa_2_i_a2_2_LC_9_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Game_Inst.r_Index_0_sqmuxa_2_i_a2_2_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__8027),
            .in2(_gnd_net_),
            .in3(N__7098),
            .lcout(\Game_Inst.N_291 ),
            .ltout(\Game_Inst.N_291_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI90L6_2_LC_9_11_5 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI90L6_2_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI90L6_2_LC_9_11_5 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \Game_Inst.r_SM_Main_RNI90L6_2_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6884),
            .in3(N__7601),
            .lcout(\Game_Inst.N_68_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Score_1_LC_9_11_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Score_1_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Score_1_LC_9_11_6 .LUT_INIT=16'b0100010101010100;
    LogicCell40 \Game_Inst.r_Score_1_LC_9_11_6  (
            .in0(N__7313),
            .in1(N__7282),
            .in2(N__7816),
            .in3(N__7859),
            .lcout(w_Score_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8259),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Score_0_LC_9_11_7 .C_ON=1'b0;
    defparam \Game_Inst.r_Score_0_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Score_0_LC_9_11_7 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \Game_Inst.r_Score_0_LC_9_11_7  (
            .in0(N__7322),
            .in1(N__7772),
            .in2(N__7283),
            .in3(N__7314),
            .lcout(w_Score_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8259),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNIERBD_0_LC_9_12_2 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNIERBD_0_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNIERBD_0_LC_9_12_2 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \Game_Inst.r_SM_Main_RNIERBD_0_LC_9_12_2  (
            .in0(N__7594),
            .in1(N__7414),
            .in2(N__7475),
            .in3(N__7700),
            .lcout(\Game_Inst.un1_r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNICE0A_0_1_LC_9_12_4 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNICE0A_0_1_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNICE0A_0_1_LC_9_12_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Game_Inst.r_SM_Main_RNICE0A_0_1_LC_9_12_4  (
            .in0(N__7595),
            .in1(N__7460),
            .in2(_gnd_net_),
            .in3(N__7413),
            .lcout(\Game_Inst.N_241 ),
            .ltout(\Game_Inst.N_241_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Score_2_LC_9_12_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Score_2_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Score_2_LC_9_12_5 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \Game_Inst.r_Score_2_LC_9_12_5  (
            .in0(N__7316),
            .in1(N__7277),
            .in2(N__7262),
            .in3(N__7259),
            .lcout(w_Score_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8264),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_9_LC_9_12_6 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_9_LC_9_12_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_9_LC_9_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_9_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7186),
            .lcout(\Game_Inst.w_LFSR_Data_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8264),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_State_e_0_LC_9_13_0 .C_ON=1'b0;
    defparam \Debounce_SW2.r_State_e_0_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_State_e_0_LC_9_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Debounce_SW2.r_State_e_0_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7156),
            .lcout(w_Switch_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8266),
            .ce(N__7136),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_State_e_0_LC_11_6_5 .C_ON=1'b0;
    defparam \Debounce_SW3.r_State_e_0_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_State_e_0_LC_11_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Debounce_SW3.r_State_e_0_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7894),
            .lcout(w_Switch_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8261),
            .ce(N__7127),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI94LD6_0_LC_11_8_1 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI94LD6_0_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI94LD6_0_LC_11_8_1 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \Game_Inst.r_SM_Main_RNI94LD6_0_LC_11_8_1  (
            .in0(N__8118),
            .in1(N__8082),
            .in2(N__7115),
            .in3(N__7980),
            .lcout(N_70),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNIBSPP6_0_LC_11_8_5 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNIBSPP6_0_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNIBSPP6_0_LC_11_8_5 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \Game_Inst.r_SM_Main_RNIBSPP6_0_LC_11_8_5  (
            .in0(N__8119),
            .in1(N__8083),
            .in2(N__7985),
            .in3(N__7937),
            .lcout(N_44),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNIC8SN6_0_LC_11_8_7 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNIC8SN6_0_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNIC8SN6_0_LC_11_8_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \Game_Inst.r_SM_Main_RNIC8SN6_0_LC_11_8_7  (
            .in0(N__8120),
            .in1(N__8084),
            .in2(N__8339),
            .in3(N__7981),
            .lcout(N_89),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_3_RNIEP6T_LC_11_9_0 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_3_RNIEP6T_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Switch_3_RNIEP6T_LC_11_9_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \Game_Inst.r_Switch_3_RNIEP6T_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__8273),
            .in2(_gnd_net_),
            .in3(N__7935),
            .lcout(\Game_Inst.N_140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_3_LC_11_9_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_3_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Switch_3_LC_11_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Switch_3_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7936),
            .lcout(\Game_Inst.r_SwitchZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8253),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNIAGNB6_0_LC_11_9_7 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNIAGNB6_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNIAGNB6_0_LC_11_9_7 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \Game_Inst.r_SM_Main_RNIAGNB6_0_LC_11_9_7  (
            .in0(N__8117),
            .in1(N__8074),
            .in2(N__8057),
            .in3(N__7979),
            .lcout(N_87),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_State_e_0_RNI8LTG1_LC_12_8_1 .C_ON=1'b0;
    defparam \Debounce_SW3.r_State_e_0_RNI8LTG1_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_State_e_0_RNI8LTG1_LC_12_8_1 .LUT_INIT=16'b1110110110100101;
    LogicCell40 \Debounce_SW3.r_State_e_0_RNI8LTG1_LC_12_8_1  (
            .in0(N__7934),
            .in1(N__7913),
            .in2(N__7901),
            .in3(N__7877),
            .lcout(\Debounce_SW3.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // State_Machine_Top
