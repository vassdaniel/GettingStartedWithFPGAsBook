-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 20 2024 18:30:00

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "Demux_Toggle_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of Demux_Toggle_TOP
entity Demux_Toggle_TOP is
port (
    o_LED_3 : out std_logic;
    o_LED_1 : out std_logic;
    i_Switch_2 : in std_logic;
    i_Clk : in std_logic;
    o_LED_4 : out std_logic;
    o_LED_2 : out std_logic;
    i_Switch_1 : in std_logic);
end Demux_Toggle_TOP;

-- Architecture of Demux_Toggle_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of Demux_Toggle_TOP is

signal \N__3212\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2655\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2566\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2524\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2456\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2449\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2395\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2388\ : std_logic;
signal \N__2385\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2353\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2340\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2332\ : std_logic;
signal \N__2331\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2295\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2284\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2254\ : std_logic;
signal \N__2251\ : std_logic;
signal \N__2248\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2233\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2212\ : std_logic;
signal \N__2211\ : std_logic;
signal \N__2208\ : std_logic;
signal \N__2205\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2190\ : std_logic;
signal \N__2187\ : std_logic;
signal \N__2184\ : std_logic;
signal \N__2181\ : std_logic;
signal \N__2178\ : std_logic;
signal \N__2175\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2167\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2163\ : std_logic;
signal \N__2160\ : std_logic;
signal \N__2157\ : std_logic;
signal \N__2154\ : std_logic;
signal \N__2147\ : std_logic;
signal \N__2144\ : std_logic;
signal \N__2141\ : std_logic;
signal \N__2138\ : std_logic;
signal \N__2135\ : std_logic;
signal \N__2132\ : std_logic;
signal \N__2131\ : std_logic;
signal \N__2128\ : std_logic;
signal \N__2125\ : std_logic;
signal \N__2122\ : std_logic;
signal \N__2119\ : std_logic;
signal \N__2114\ : std_logic;
signal \N__2111\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2109\ : std_logic;
signal \N__2106\ : std_logic;
signal \N__2105\ : std_logic;
signal \N__2104\ : std_logic;
signal \N__2101\ : std_logic;
signal \N__2100\ : std_logic;
signal \N__2097\ : std_logic;
signal \N__2094\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2087\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2085\ : std_logic;
signal \N__2078\ : std_logic;
signal \N__2073\ : std_logic;
signal \N__2070\ : std_logic;
signal \N__2065\ : std_logic;
signal \N__2062\ : std_logic;
signal \N__2051\ : std_logic;
signal \N__2050\ : std_logic;
signal \N__2049\ : std_logic;
signal \N__2048\ : std_logic;
signal \N__2045\ : std_logic;
signal \N__2044\ : std_logic;
signal \N__2043\ : std_logic;
signal \N__2042\ : std_logic;
signal \N__2041\ : std_logic;
signal \N__2038\ : std_logic;
signal \N__2035\ : std_logic;
signal \N__2028\ : std_logic;
signal \N__2025\ : std_logic;
signal \N__2020\ : std_logic;
signal \N__2009\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2003\ : std_logic;
signal \N__2002\ : std_logic;
signal \N__1999\ : std_logic;
signal \N__1996\ : std_logic;
signal \N__1991\ : std_logic;
signal \N__1990\ : std_logic;
signal \N__1987\ : std_logic;
signal \N__1984\ : std_logic;
signal \N__1979\ : std_logic;
signal \N__1978\ : std_logic;
signal \N__1977\ : std_logic;
signal \N__1972\ : std_logic;
signal \N__1969\ : std_logic;
signal \N__1964\ : std_logic;
signal \N__1961\ : std_logic;
signal \N__1958\ : std_logic;
signal \N__1955\ : std_logic;
signal \N__1952\ : std_logic;
signal \N__1951\ : std_logic;
signal \N__1948\ : std_logic;
signal \N__1945\ : std_logic;
signal \N__1940\ : std_logic;
signal \N__1937\ : std_logic;
signal \N__1934\ : std_logic;
signal \N__1933\ : std_logic;
signal \N__1930\ : std_logic;
signal \N__1927\ : std_logic;
signal \N__1924\ : std_logic;
signal \N__1921\ : std_logic;
signal \N__1916\ : std_logic;
signal \N__1915\ : std_logic;
signal \N__1912\ : std_logic;
signal \N__1909\ : std_logic;
signal \N__1904\ : std_logic;
signal \N__1901\ : std_logic;
signal \N__1898\ : std_logic;
signal \N__1895\ : std_logic;
signal \N__1894\ : std_logic;
signal \N__1891\ : std_logic;
signal \N__1888\ : std_logic;
signal \N__1883\ : std_logic;
signal \N__1882\ : std_logic;
signal \N__1879\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1871\ : std_logic;
signal \N__1870\ : std_logic;
signal \N__1867\ : std_logic;
signal \N__1864\ : std_logic;
signal \N__1859\ : std_logic;
signal \N__1858\ : std_logic;
signal \N__1857\ : std_logic;
signal \N__1856\ : std_logic;
signal \N__1853\ : std_logic;
signal \N__1848\ : std_logic;
signal \N__1845\ : std_logic;
signal \N__1842\ : std_logic;
signal \N__1835\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1829\ : std_logic;
signal \N__1826\ : std_logic;
signal \N__1823\ : std_logic;
signal \N__1820\ : std_logic;
signal \N__1817\ : std_logic;
signal \N__1814\ : std_logic;
signal \N__1811\ : std_logic;
signal \N__1808\ : std_logic;
signal \N__1805\ : std_logic;
signal \N__1802\ : std_logic;
signal \N__1801\ : std_logic;
signal \N__1800\ : std_logic;
signal \N__1799\ : std_logic;
signal \N__1790\ : std_logic;
signal \N__1787\ : std_logic;
signal \N__1784\ : std_logic;
signal \N__1781\ : std_logic;
signal \N__1780\ : std_logic;
signal \N__1777\ : std_logic;
signal \N__1774\ : std_logic;
signal \N__1769\ : std_logic;
signal \N__1768\ : std_logic;
signal \N__1765\ : std_logic;
signal \N__1762\ : std_logic;
signal \N__1757\ : std_logic;
signal \N__1754\ : std_logic;
signal \N__1753\ : std_logic;
signal \N__1750\ : std_logic;
signal \N__1747\ : std_logic;
signal \N__1742\ : std_logic;
signal \N__1741\ : std_logic;
signal \N__1738\ : std_logic;
signal \N__1735\ : std_logic;
signal \N__1730\ : std_logic;
signal \N__1727\ : std_logic;
signal \N__1724\ : std_logic;
signal \N__1723\ : std_logic;
signal \N__1720\ : std_logic;
signal \N__1717\ : std_logic;
signal \N__1714\ : std_logic;
signal \N__1709\ : std_logic;
signal \N__1708\ : std_logic;
signal \N__1705\ : std_logic;
signal \N__1702\ : std_logic;
signal \N__1697\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1693\ : std_logic;
signal \N__1690\ : std_logic;
signal \N__1685\ : std_logic;
signal \N__1684\ : std_logic;
signal \N__1681\ : std_logic;
signal \N__1678\ : std_logic;
signal \N__1673\ : std_logic;
signal \N__1670\ : std_logic;
signal \N__1667\ : std_logic;
signal \N__1664\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1658\ : std_logic;
signal \N__1655\ : std_logic;
signal \N__1652\ : std_logic;
signal \N__1649\ : std_logic;
signal \N__1646\ : std_logic;
signal \N__1643\ : std_logic;
signal \N__1640\ : std_logic;
signal \N__1637\ : std_logic;
signal \N__1634\ : std_logic;
signal \N__1633\ : std_logic;
signal \N__1628\ : std_logic;
signal \N__1625\ : std_logic;
signal \N__1624\ : std_logic;
signal \N__1619\ : std_logic;
signal \N__1616\ : std_logic;
signal \N__1613\ : std_logic;
signal \N__1612\ : std_logic;
signal \N__1607\ : std_logic;
signal \N__1604\ : std_logic;
signal \N__1603\ : std_logic;
signal \N__1598\ : std_logic;
signal \N__1595\ : std_logic;
signal \N__1594\ : std_logic;
signal \N__1593\ : std_logic;
signal \N__1592\ : std_logic;
signal \N__1589\ : std_logic;
signal \N__1582\ : std_logic;
signal \N__1577\ : std_logic;
signal \N__1576\ : std_logic;
signal \N__1573\ : std_logic;
signal \N__1570\ : std_logic;
signal \N__1569\ : std_logic;
signal \N__1566\ : std_logic;
signal \N__1561\ : std_logic;
signal \N__1556\ : std_logic;
signal \N__1555\ : std_logic;
signal \N__1552\ : std_logic;
signal \N__1549\ : std_logic;
signal \N__1544\ : std_logic;
signal \N__1541\ : std_logic;
signal \N__1540\ : std_logic;
signal \N__1537\ : std_logic;
signal \N__1534\ : std_logic;
signal \N__1531\ : std_logic;
signal \N__1526\ : std_logic;
signal \N__1523\ : std_logic;
signal \N__1522\ : std_logic;
signal \N__1519\ : std_logic;
signal \N__1516\ : std_logic;
signal \N__1511\ : std_logic;
signal \N__1508\ : std_logic;
signal \N__1505\ : std_logic;
signal \N__1502\ : std_logic;
signal \N__1499\ : std_logic;
signal \N__1496\ : std_logic;
signal \N__1493\ : std_logic;
signal \N__1490\ : std_logic;
signal \N__1487\ : std_logic;
signal \N__1484\ : std_logic;
signal \N__1481\ : std_logic;
signal \N__1478\ : std_logic;
signal \N__1475\ : std_logic;
signal \N__1472\ : std_logic;
signal \N__1469\ : std_logic;
signal \N__1466\ : std_logic;
signal \N__1463\ : std_logic;
signal \N__1460\ : std_logic;
signal \N__1457\ : std_logic;
signal \N__1454\ : std_logic;
signal \N__1451\ : std_logic;
signal \N__1448\ : std_logic;
signal \N__1445\ : std_logic;
signal \N__1442\ : std_logic;
signal \N__1439\ : std_logic;
signal \N__1436\ : std_logic;
signal \N__1433\ : std_logic;
signal \N__1430\ : std_logic;
signal \N__1427\ : std_logic;
signal \N__1424\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \Debounce_Sw1.un9_r_count_10_cascade_\ : std_logic;
signal \Debounce_Sw1.un1_r_Count_1lt11_0_cascade_\ : std_logic;
signal \Debounce_Sw1.un1_r_Count_1lto11_1\ : std_logic;
signal \Debounce_Sw1.un1_r_Count_1lt17_cascade_\ : std_logic;
signal \Debounce_Sw1.un1_r_Count_1lto17_2\ : std_logic;
signal \Debounce_Sw1.r_count15_i\ : std_logic;
signal \bfn_4_7_0_\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_1\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_2\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_3\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_4\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_5\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_6\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_7\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_8\ : std_logic;
signal \bfn_4_8_0_\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_9\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_10\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_11\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_12\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_13\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_14\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_15\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_16\ : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_17\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_18\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_19\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_20\ : std_logic;
signal \Count_And_Toggle.un2_r_counter_cry_21\ : std_logic;
signal \Count_And_Toggle.r_Counter_RNO_0Z0Z_22_cascade_\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_17\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_22\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_21\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_20\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_0\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_1\ : std_logic;
signal \bfn_5_5_0_\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_2\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_1\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_3\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_2\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_4\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_3\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_5\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_4\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_5\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_6\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_7\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_8\ : std_logic;
signal \bfn_5_6_0_\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_9\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_10\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_11\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_12\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_13\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_14\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_15\ : std_logic;
signal \Debounce_Sw1.un2_r_count_cry_16\ : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal \Debounce_Sw1.r_count15_i_g\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_12\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_10\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_13\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_7\ : std_logic;
signal \Count_And_Toggle.r_Counter_RNO_0Z0Z_8\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_8\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_5\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_4\ : std_logic;
signal \Count_And_Toggle.r_Counter_RNO_0Z0Z_11\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_3\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_2\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_1\ : std_logic;
signal \Count_And_Toggle.r_Counter_RNO_0Z0Z_6\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_6\ : std_logic;
signal \Count_And_Toggle.r_Counter_RNO_0Z0Z_19\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_19\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_11\ : std_logic;
signal \Count_And_Toggle.un4_i_enable_15_cascade_\ : std_logic;
signal \Count_And_Toggle.r_Counter_RNO_0Z0Z_18\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_18\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_15\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_16\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_0\ : std_logic;
signal \Count_And_Toggle.un4_i_enable_14\ : std_logic;
signal \Count_And_Toggle.un4_i_enable_12\ : std_logic;
signal \Count_And_Toggle.un4_i_enable_11_cascade_\ : std_logic;
signal \Count_And_Toggle.un4_i_enable_13\ : std_logic;
signal \Count_And_Toggle.un4_i_enable_20_cascade_\ : std_logic;
signal \Count_And_Toggle.r_Counter_RNO_0Z0Z_14\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_14\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_8\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_6\ : std_logic;
signal \Debounce_Sw1.un9_r_count_9\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_12\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_14\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_15\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_7\ : std_logic;
signal \Debounce_Sw1.un9_r_count_10\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_9\ : std_logic;
signal \Debounce_Sw1.un9_r_count_5_cascade_\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_10\ : std_logic;
signal \Debounce_Sw1.un9_r_count_9_0\ : std_logic;
signal \i_Switch_1_c\ : std_logic;
signal \Debounce_Sw1.un9_r_count_10_0_cascade_\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_16\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_13\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_17\ : std_logic;
signal \Debounce_Sw1.r_CountZ0Z_11\ : std_logic;
signal \Debounce_Sw1.un9_r_count_6\ : std_logic;
signal \Count_And_Toggle.r_Counter_RNO_0Z0Z_9\ : std_logic;
signal \Count_And_Toggle.r_CounterZ0Z_9\ : std_logic;
signal \Count_And_Toggle.un4_i_enable_16\ : std_logic;
signal \Count_And_Toggle.un4_i_enable_15\ : std_logic;
signal \Count_And_Toggle.un4_i_enable_20\ : std_logic;
signal \Debounce_Sw2.un9_r_count_10_cascade_\ : std_logic;
signal \Debounce_Sw2.N_23_cascade_\ : std_logic;
signal \i_Switch_2_c\ : std_logic;
signal \Debounce_Sw2.N_16_cascade_\ : std_logic;
signal \Debounce_Sw2.N_9\ : std_logic;
signal \Debounce_Sw2.un9_r_count_10\ : std_logic;
signal \Debounce_Sw2.r_State_e_0_RNOZ0\ : std_logic;
signal \Debounce_Sw2.N_10\ : std_logic;
signal \Debounce_Sw2.un9_r_count_0_a3_2\ : std_logic;
signal \Debounce_Sw2.N_22_3\ : std_logic;
signal \Debounce_Sw2.N_13\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_0\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_1\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_2\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_1\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_3\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_2\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_4\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_3\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_5\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_4\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_6\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_5\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_7\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_6\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_8\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_7\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_8\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_9\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_10\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_9\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_11\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_10\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_12\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_11\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_13\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_12\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_14\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_13\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_15\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_14\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_16\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_15\ : std_logic;
signal \Debounce_Sw2.un2_r_count_cry_16\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \Debounce_Sw2.r_CountZ0Z_17\ : std_logic;
signal \i_Clk_c_g\ : std_logic;
signal \Debounce_Sw2.N_9_g\ : std_logic;
signal \o_LED_2_c\ : std_logic;
signal \o_LED_3_c\ : std_logic;
signal \o_LED_1_c\ : std_logic;
signal \w_Switch_1\ : std_logic;
signal \w_Toggle\ : std_logic;
signal \w_Switch_2\ : std_logic;
signal \o_LED_4_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \i_Clk_wire\ : std_logic;
signal \o_LED_1_wire\ : std_logic;
signal \i_Switch_1_wire\ : std_logic;
signal \o_LED_2_wire\ : std_logic;
signal \i_Switch_2_wire\ : std_logic;
signal \o_LED_3_wire\ : std_logic;
signal \o_LED_4_wire\ : std_logic;

begin
    \i_Clk_wire\ <= i_Clk;
    o_LED_1 <= \o_LED_1_wire\;
    \i_Switch_1_wire\ <= i_Switch_1;
    o_LED_2 <= \o_LED_2_wire\;
    \i_Switch_2_wire\ <= i_Switch_2;
    o_LED_3 <= \o_LED_3_wire\;
    o_LED_4 <= \o_LED_4_wire\;

    \i_Clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__3210\,
            GLOBALBUFFEROUTPUT => \i_Clk_c_g\
        );

    \i_Clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3212\,
            DIN => \N__3211\,
            DOUT => \N__3210\,
            PACKAGEPIN => \i_Clk_wire\
        );

    \i_Clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3212\,
            PADOUT => \N__3211\,
            PADIN => \N__3210\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3201\,
            DIN => \N__3200\,
            DOUT => \N__3199\,
            PACKAGEPIN => \o_LED_1_wire\
        );

    \o_LED_1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3201\,
            PADOUT => \N__3200\,
            PADIN => \N__3199\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2999\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_Switch_1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3192\,
            DIN => \N__3191\,
            DOUT => \N__3190\,
            PACKAGEPIN => \i_Switch_1_wire\
        );

    \i_Switch_1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3192\,
            PADOUT => \N__3191\,
            PADIN => \N__3190\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \i_Switch_1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3183\,
            DIN => \N__3182\,
            DOUT => \N__3181\,
            PACKAGEPIN => \o_LED_2_wire\
        );

    \o_LED_2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3183\,
            PADOUT => \N__3182\,
            PADIN => \N__3181\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3011\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_Switch_2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3174\,
            DIN => \N__3173\,
            DOUT => \N__3172\,
            PACKAGEPIN => \i_Switch_2_wire\
        );

    \i_Switch_2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3174\,
            PADOUT => \N__3173\,
            PADIN => \N__3172\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \i_Switch_2_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3165\,
            DIN => \N__3164\,
            DOUT => \N__3163\,
            PACKAGEPIN => \o_LED_3_wire\
        );

    \o_LED_3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3165\,
            PADOUT => \N__3164\,
            PADIN => \N__3163\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3005\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3156\,
            DIN => \N__3155\,
            DOUT => \N__3154\,
            PACKAGEPIN => \o_LED_4_wire\
        );

    \o_LED_4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3156\,
            PADOUT => \N__3155\,
            PADIN => \N__3154\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2882\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__696\ : InMux
    port map (
            O => \N__3137\,
            I => \N__3133\
        );

    \I__695\ : InMux
    port map (
            O => \N__3136\,
            I => \N__3130\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3133\,
            I => \Debounce_Sw2.r_CountZ0Z_15\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3130\,
            I => \Debounce_Sw2.r_CountZ0Z_15\
        );

    \I__692\ : InMux
    port map (
            O => \N__3125\,
            I => \Debounce_Sw2.un2_r_count_cry_14\
        );

    \I__691\ : InMux
    port map (
            O => \N__3122\,
            I => \N__3118\
        );

    \I__690\ : InMux
    port map (
            O => \N__3121\,
            I => \N__3115\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3118\,
            I => \Debounce_Sw2.r_CountZ0Z_16\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3115\,
            I => \Debounce_Sw2.r_CountZ0Z_16\
        );

    \I__687\ : InMux
    port map (
            O => \N__3110\,
            I => \Debounce_Sw2.un2_r_count_cry_15\
        );

    \I__686\ : InMux
    port map (
            O => \N__3107\,
            I => \bfn_8_11_0_\
        );

    \I__685\ : CascadeMux
    port map (
            O => \N__3104\,
            I => \N__3101\
        );

    \I__684\ : InMux
    port map (
            O => \N__3101\,
            I => \N__3097\
        );

    \I__683\ : InMux
    port map (
            O => \N__3100\,
            I => \N__3094\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__3097\,
            I => \N__3091\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3094\,
            I => \Debounce_Sw2.r_CountZ0Z_17\
        );

    \I__680\ : Odrv4
    port map (
            O => \N__3091\,
            I => \Debounce_Sw2.r_CountZ0Z_17\
        );

    \I__679\ : ClkMux
    port map (
            O => \N__3086\,
            I => \N__3035\
        );

    \I__678\ : ClkMux
    port map (
            O => \N__3085\,
            I => \N__3035\
        );

    \I__677\ : ClkMux
    port map (
            O => \N__3084\,
            I => \N__3035\
        );

    \I__676\ : ClkMux
    port map (
            O => \N__3083\,
            I => \N__3035\
        );

    \I__675\ : ClkMux
    port map (
            O => \N__3082\,
            I => \N__3035\
        );

    \I__674\ : ClkMux
    port map (
            O => \N__3081\,
            I => \N__3035\
        );

    \I__673\ : ClkMux
    port map (
            O => \N__3080\,
            I => \N__3035\
        );

    \I__672\ : ClkMux
    port map (
            O => \N__3079\,
            I => \N__3035\
        );

    \I__671\ : ClkMux
    port map (
            O => \N__3078\,
            I => \N__3035\
        );

    \I__670\ : ClkMux
    port map (
            O => \N__3077\,
            I => \N__3035\
        );

    \I__669\ : ClkMux
    port map (
            O => \N__3076\,
            I => \N__3035\
        );

    \I__668\ : ClkMux
    port map (
            O => \N__3075\,
            I => \N__3035\
        );

    \I__667\ : ClkMux
    port map (
            O => \N__3074\,
            I => \N__3035\
        );

    \I__666\ : ClkMux
    port map (
            O => \N__3073\,
            I => \N__3035\
        );

    \I__665\ : ClkMux
    port map (
            O => \N__3072\,
            I => \N__3035\
        );

    \I__664\ : ClkMux
    port map (
            O => \N__3071\,
            I => \N__3035\
        );

    \I__663\ : ClkMux
    port map (
            O => \N__3070\,
            I => \N__3035\
        );

    \I__662\ : GlobalMux
    port map (
            O => \N__3035\,
            I => \N__3032\
        );

    \I__661\ : gio2CtrlBuf
    port map (
            O => \N__3032\,
            I => \i_Clk_c_g\
        );

    \I__660\ : SRMux
    port map (
            O => \N__3029\,
            I => \N__3017\
        );

    \I__659\ : SRMux
    port map (
            O => \N__3028\,
            I => \N__3017\
        );

    \I__658\ : SRMux
    port map (
            O => \N__3027\,
            I => \N__3017\
        );

    \I__657\ : SRMux
    port map (
            O => \N__3026\,
            I => \N__3017\
        );

    \I__656\ : GlobalMux
    port map (
            O => \N__3017\,
            I => \N__3014\
        );

    \I__655\ : gio2CtrlBuf
    port map (
            O => \N__3014\,
            I => \Debounce_Sw2.N_9_g\
        );

    \I__654\ : IoInMux
    port map (
            O => \N__3011\,
            I => \N__3008\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3008\,
            I => \o_LED_2_c\
        );

    \I__652\ : IoInMux
    port map (
            O => \N__3005\,
            I => \N__3002\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3002\,
            I => \o_LED_3_c\
        );

    \I__650\ : IoInMux
    port map (
            O => \N__2999\,
            I => \N__2996\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__2996\,
            I => \o_LED_1_c\
        );

    \I__648\ : InMux
    port map (
            O => \N__2993\,
            I => \N__2987\
        );

    \I__647\ : InMux
    port map (
            O => \N__2992\,
            I => \N__2980\
        );

    \I__646\ : InMux
    port map (
            O => \N__2991\,
            I => \N__2980\
        );

    \I__645\ : InMux
    port map (
            O => \N__2990\,
            I => \N__2980\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__2987\,
            I => \N__2975\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__2980\,
            I => \N__2975\
        );

    \I__642\ : Span4Mux_v
    port map (
            O => \N__2975\,
            I => \N__2970\
        );

    \I__641\ : InMux
    port map (
            O => \N__2974\,
            I => \N__2967\
        );

    \I__640\ : InMux
    port map (
            O => \N__2973\,
            I => \N__2964\
        );

    \I__639\ : Span4Mux_h
    port map (
            O => \N__2970\,
            I => \N__2959\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__2967\,
            I => \N__2959\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__2964\,
            I => \w_Switch_1\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__2959\,
            I => \w_Switch_1\
        );

    \I__635\ : InMux
    port map (
            O => \N__2954\,
            I => \N__2944\
        );

    \I__634\ : InMux
    port map (
            O => \N__2953\,
            I => \N__2944\
        );

    \I__633\ : InMux
    port map (
            O => \N__2952\,
            I => \N__2944\
        );

    \I__632\ : InMux
    port map (
            O => \N__2951\,
            I => \N__2941\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__2944\,
            I => \N__2936\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__2941\,
            I => \N__2936\
        );

    \I__629\ : Span4Mux_v
    port map (
            O => \N__2936\,
            I => \N__2932\
        );

    \I__628\ : CascadeMux
    port map (
            O => \N__2935\,
            I => \N__2929\
        );

    \I__627\ : Span4Mux_h
    port map (
            O => \N__2932\,
            I => \N__2926\
        );

    \I__626\ : InMux
    port map (
            O => \N__2929\,
            I => \N__2923\
        );

    \I__625\ : Odrv4
    port map (
            O => \N__2926\,
            I => \w_Toggle\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__2923\,
            I => \w_Toggle\
        );

    \I__623\ : CascadeMux
    port map (
            O => \N__2918\,
            I => \N__2914\
        );

    \I__622\ : InMux
    port map (
            O => \N__2917\,
            I => \N__2905\
        );

    \I__621\ : InMux
    port map (
            O => \N__2914\,
            I => \N__2905\
        );

    \I__620\ : InMux
    port map (
            O => \N__2913\,
            I => \N__2905\
        );

    \I__619\ : InMux
    port map (
            O => \N__2912\,
            I => \N__2902\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__2905\,
            I => \N__2897\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__2902\,
            I => \N__2897\
        );

    \I__616\ : Span4Mux_v
    port map (
            O => \N__2897\,
            I => \N__2894\
        );

    \I__615\ : Span4Mux_h
    port map (
            O => \N__2894\,
            I => \N__2890\
        );

    \I__614\ : InMux
    port map (
            O => \N__2893\,
            I => \N__2887\
        );

    \I__613\ : Odrv4
    port map (
            O => \N__2890\,
            I => \w_Switch_2\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__2887\,
            I => \w_Switch_2\
        );

    \I__611\ : IoInMux
    port map (
            O => \N__2882\,
            I => \N__2879\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__2879\,
            I => \o_LED_4_c\
        );

    \I__609\ : InMux
    port map (
            O => \N__2876\,
            I => \N__2872\
        );

    \I__608\ : InMux
    port map (
            O => \N__2875\,
            I => \N__2869\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__2872\,
            I => \Debounce_Sw2.r_CountZ0Z_6\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__2869\,
            I => \Debounce_Sw2.r_CountZ0Z_6\
        );

    \I__605\ : InMux
    port map (
            O => \N__2864\,
            I => \Debounce_Sw2.un2_r_count_cry_5\
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__2861\,
            I => \N__2857\
        );

    \I__603\ : InMux
    port map (
            O => \N__2860\,
            I => \N__2853\
        );

    \I__602\ : InMux
    port map (
            O => \N__2857\,
            I => \N__2850\
        );

    \I__601\ : InMux
    port map (
            O => \N__2856\,
            I => \N__2847\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__2853\,
            I => \Debounce_Sw2.r_CountZ0Z_7\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__2850\,
            I => \Debounce_Sw2.r_CountZ0Z_7\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__2847\,
            I => \Debounce_Sw2.r_CountZ0Z_7\
        );

    \I__597\ : InMux
    port map (
            O => \N__2840\,
            I => \Debounce_Sw2.un2_r_count_cry_6\
        );

    \I__596\ : InMux
    port map (
            O => \N__2837\,
            I => \N__2833\
        );

    \I__595\ : InMux
    port map (
            O => \N__2836\,
            I => \N__2830\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__2833\,
            I => \Debounce_Sw2.r_CountZ0Z_8\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__2830\,
            I => \Debounce_Sw2.r_CountZ0Z_8\
        );

    \I__592\ : InMux
    port map (
            O => \N__2825\,
            I => \Debounce_Sw2.un2_r_count_cry_7\
        );

    \I__591\ : InMux
    port map (
            O => \N__2822\,
            I => \N__2818\
        );

    \I__590\ : InMux
    port map (
            O => \N__2821\,
            I => \N__2815\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__2818\,
            I => \Debounce_Sw2.r_CountZ0Z_9\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__2815\,
            I => \Debounce_Sw2.r_CountZ0Z_9\
        );

    \I__587\ : InMux
    port map (
            O => \N__2810\,
            I => \bfn_8_10_0_\
        );

    \I__586\ : InMux
    port map (
            O => \N__2807\,
            I => \N__2803\
        );

    \I__585\ : InMux
    port map (
            O => \N__2806\,
            I => \N__2800\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__2803\,
            I => \Debounce_Sw2.r_CountZ0Z_10\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__2800\,
            I => \Debounce_Sw2.r_CountZ0Z_10\
        );

    \I__582\ : InMux
    port map (
            O => \N__2795\,
            I => \Debounce_Sw2.un2_r_count_cry_9\
        );

    \I__581\ : CascadeMux
    port map (
            O => \N__2792\,
            I => \N__2788\
        );

    \I__580\ : InMux
    port map (
            O => \N__2791\,
            I => \N__2785\
        );

    \I__579\ : InMux
    port map (
            O => \N__2788\,
            I => \N__2782\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__2785\,
            I => \Debounce_Sw2.r_CountZ0Z_11\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__2782\,
            I => \Debounce_Sw2.r_CountZ0Z_11\
        );

    \I__576\ : InMux
    port map (
            O => \N__2777\,
            I => \Debounce_Sw2.un2_r_count_cry_10\
        );

    \I__575\ : InMux
    port map (
            O => \N__2774\,
            I => \N__2769\
        );

    \I__574\ : InMux
    port map (
            O => \N__2773\,
            I => \N__2764\
        );

    \I__573\ : InMux
    port map (
            O => \N__2772\,
            I => \N__2764\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__2769\,
            I => \Debounce_Sw2.r_CountZ0Z_12\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__2764\,
            I => \Debounce_Sw2.r_CountZ0Z_12\
        );

    \I__570\ : InMux
    port map (
            O => \N__2759\,
            I => \Debounce_Sw2.un2_r_count_cry_11\
        );

    \I__569\ : InMux
    port map (
            O => \N__2756\,
            I => \N__2751\
        );

    \I__568\ : InMux
    port map (
            O => \N__2755\,
            I => \N__2748\
        );

    \I__567\ : InMux
    port map (
            O => \N__2754\,
            I => \N__2745\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__2751\,
            I => \Debounce_Sw2.r_CountZ0Z_13\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__2748\,
            I => \Debounce_Sw2.r_CountZ0Z_13\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__2745\,
            I => \Debounce_Sw2.r_CountZ0Z_13\
        );

    \I__563\ : InMux
    port map (
            O => \N__2738\,
            I => \Debounce_Sw2.un2_r_count_cry_12\
        );

    \I__562\ : InMux
    port map (
            O => \N__2735\,
            I => \N__2731\
        );

    \I__561\ : InMux
    port map (
            O => \N__2734\,
            I => \N__2728\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__2731\,
            I => \Debounce_Sw2.r_CountZ0Z_14\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__2728\,
            I => \Debounce_Sw2.r_CountZ0Z_14\
        );

    \I__558\ : InMux
    port map (
            O => \N__2723\,
            I => \Debounce_Sw2.un2_r_count_cry_13\
        );

    \I__557\ : InMux
    port map (
            O => \N__2720\,
            I => \N__2716\
        );

    \I__556\ : InMux
    port map (
            O => \N__2719\,
            I => \N__2713\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__2716\,
            I => \Debounce_Sw2.N_10\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__2713\,
            I => \Debounce_Sw2.N_10\
        );

    \I__553\ : InMux
    port map (
            O => \N__2708\,
            I => \N__2705\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__2705\,
            I => \Debounce_Sw2.un9_r_count_0_a3_2\
        );

    \I__551\ : InMux
    port map (
            O => \N__2702\,
            I => \N__2696\
        );

    \I__550\ : InMux
    port map (
            O => \N__2701\,
            I => \N__2696\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__2696\,
            I => \Debounce_Sw2.N_22_3\
        );

    \I__548\ : InMux
    port map (
            O => \N__2693\,
            I => \N__2687\
        );

    \I__547\ : InMux
    port map (
            O => \N__2692\,
            I => \N__2687\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__2687\,
            I => \Debounce_Sw2.N_13\
        );

    \I__545\ : InMux
    port map (
            O => \N__2684\,
            I => \N__2676\
        );

    \I__544\ : InMux
    port map (
            O => \N__2683\,
            I => \N__2676\
        );

    \I__543\ : InMux
    port map (
            O => \N__2682\,
            I => \N__2673\
        );

    \I__542\ : InMux
    port map (
            O => \N__2681\,
            I => \N__2670\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__2676\,
            I => \Debounce_Sw2.r_CountZ0Z_0\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__2673\,
            I => \Debounce_Sw2.r_CountZ0Z_0\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__2670\,
            I => \Debounce_Sw2.r_CountZ0Z_0\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__2663\,
            I => \N__2659\
        );

    \I__537\ : InMux
    port map (
            O => \N__2662\,
            I => \N__2655\
        );

    \I__536\ : InMux
    port map (
            O => \N__2659\,
            I => \N__2652\
        );

    \I__535\ : InMux
    port map (
            O => \N__2658\,
            I => \N__2649\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__2655\,
            I => \Debounce_Sw2.r_CountZ0Z_1\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__2652\,
            I => \Debounce_Sw2.r_CountZ0Z_1\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__2649\,
            I => \Debounce_Sw2.r_CountZ0Z_1\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__2642\,
            I => \N__2639\
        );

    \I__530\ : InMux
    port map (
            O => \N__2639\,
            I => \N__2635\
        );

    \I__529\ : InMux
    port map (
            O => \N__2638\,
            I => \N__2632\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__2635\,
            I => \N__2629\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__2632\,
            I => \Debounce_Sw2.r_CountZ0Z_2\
        );

    \I__526\ : Odrv4
    port map (
            O => \N__2629\,
            I => \Debounce_Sw2.r_CountZ0Z_2\
        );

    \I__525\ : InMux
    port map (
            O => \N__2624\,
            I => \Debounce_Sw2.un2_r_count_cry_1\
        );

    \I__524\ : InMux
    port map (
            O => \N__2621\,
            I => \N__2617\
        );

    \I__523\ : InMux
    port map (
            O => \N__2620\,
            I => \N__2614\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__2617\,
            I => \Debounce_Sw2.r_CountZ0Z_3\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__2614\,
            I => \Debounce_Sw2.r_CountZ0Z_3\
        );

    \I__520\ : InMux
    port map (
            O => \N__2609\,
            I => \Debounce_Sw2.un2_r_count_cry_2\
        );

    \I__519\ : InMux
    port map (
            O => \N__2606\,
            I => \N__2602\
        );

    \I__518\ : InMux
    port map (
            O => \N__2605\,
            I => \N__2599\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__2602\,
            I => \Debounce_Sw2.r_CountZ0Z_4\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__2599\,
            I => \Debounce_Sw2.r_CountZ0Z_4\
        );

    \I__515\ : InMux
    port map (
            O => \N__2594\,
            I => \Debounce_Sw2.un2_r_count_cry_3\
        );

    \I__514\ : InMux
    port map (
            O => \N__2591\,
            I => \N__2587\
        );

    \I__513\ : InMux
    port map (
            O => \N__2590\,
            I => \N__2584\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__2587\,
            I => \N__2581\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__2584\,
            I => \Debounce_Sw2.r_CountZ0Z_5\
        );

    \I__510\ : Odrv4
    port map (
            O => \N__2581\,
            I => \Debounce_Sw2.r_CountZ0Z_5\
        );

    \I__509\ : InMux
    port map (
            O => \N__2576\,
            I => \Debounce_Sw2.un2_r_count_cry_4\
        );

    \I__508\ : InMux
    port map (
            O => \N__2573\,
            I => \N__2563\
        );

    \I__507\ : InMux
    port map (
            O => \N__2572\,
            I => \N__2560\
        );

    \I__506\ : InMux
    port map (
            O => \N__2571\,
            I => \N__2553\
        );

    \I__505\ : InMux
    port map (
            O => \N__2570\,
            I => \N__2553\
        );

    \I__504\ : InMux
    port map (
            O => \N__2569\,
            I => \N__2553\
        );

    \I__503\ : InMux
    port map (
            O => \N__2568\,
            I => \N__2550\
        );

    \I__502\ : InMux
    port map (
            O => \N__2567\,
            I => \N__2545\
        );

    \I__501\ : InMux
    port map (
            O => \N__2566\,
            I => \N__2545\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__2563\,
            I => \Count_And_Toggle.un4_i_enable_20\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__2560\,
            I => \Count_And_Toggle.un4_i_enable_20\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__2553\,
            I => \Count_And_Toggle.un4_i_enable_20\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__2550\,
            I => \Count_And_Toggle.un4_i_enable_20\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__2545\,
            I => \Count_And_Toggle.un4_i_enable_20\
        );

    \I__495\ : CascadeMux
    port map (
            O => \N__2534\,
            I => \Debounce_Sw2.un9_r_count_10_cascade_\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__2531\,
            I => \Debounce_Sw2.N_23_cascade_\
        );

    \I__493\ : InMux
    port map (
            O => \N__2528\,
            I => \N__2525\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__2525\,
            I => \N__2521\
        );

    \I__491\ : InMux
    port map (
            O => \N__2524\,
            I => \N__2518\
        );

    \I__490\ : Span4Mux_v
    port map (
            O => \N__2521\,
            I => \N__2515\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__2518\,
            I => \N__2512\
        );

    \I__488\ : Span4Mux_h
    port map (
            O => \N__2515\,
            I => \N__2509\
        );

    \I__487\ : Span12Mux_v
    port map (
            O => \N__2512\,
            I => \N__2506\
        );

    \I__486\ : Span4Mux_v
    port map (
            O => \N__2509\,
            I => \N__2503\
        );

    \I__485\ : Odrv12
    port map (
            O => \N__2506\,
            I => \i_Switch_2_c\
        );

    \I__484\ : Odrv4
    port map (
            O => \N__2503\,
            I => \i_Switch_2_c\
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__2498\,
            I => \Debounce_Sw2.N_16_cascade_\
        );

    \I__482\ : IoInMux
    port map (
            O => \N__2495\,
            I => \N__2492\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2492\,
            I => \N__2489\
        );

    \I__480\ : Span12Mux_s7_v
    port map (
            O => \N__2489\,
            I => \N__2486\
        );

    \I__479\ : Odrv12
    port map (
            O => \N__2486\,
            I => \Debounce_Sw2.N_9\
        );

    \I__478\ : CascadeMux
    port map (
            O => \N__2483\,
            I => \N__2480\
        );

    \I__477\ : InMux
    port map (
            O => \N__2480\,
            I => \N__2477\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__2477\,
            I => \Debounce_Sw2.un9_r_count_10\
        );

    \I__475\ : CEMux
    port map (
            O => \N__2474\,
            I => \N__2471\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__2471\,
            I => \N__2468\
        );

    \I__473\ : Odrv4
    port map (
            O => \N__2468\,
            I => \Debounce_Sw2.r_State_e_0_RNOZ0\
        );

    \I__472\ : CascadeMux
    port map (
            O => \N__2465\,
            I => \Count_And_Toggle.un4_i_enable_20_cascade_\
        );

    \I__471\ : InMux
    port map (
            O => \N__2462\,
            I => \N__2459\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__2459\,
            I => \Count_And_Toggle.r_Counter_RNO_0Z0Z_14\
        );

    \I__469\ : InMux
    port map (
            O => \N__2456\,
            I => \N__2452\
        );

    \I__468\ : InMux
    port map (
            O => \N__2455\,
            I => \N__2449\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__2452\,
            I => \Count_And_Toggle.r_CounterZ0Z_14\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__2449\,
            I => \Count_And_Toggle.r_CounterZ0Z_14\
        );

    \I__465\ : InMux
    port map (
            O => \N__2444\,
            I => \N__2439\
        );

    \I__464\ : InMux
    port map (
            O => \N__2443\,
            I => \N__2436\
        );

    \I__463\ : InMux
    port map (
            O => \N__2442\,
            I => \N__2433\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2439\,
            I => \Debounce_Sw1.r_CountZ0Z_8\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__2436\,
            I => \Debounce_Sw1.r_CountZ0Z_8\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__2433\,
            I => \Debounce_Sw1.r_CountZ0Z_8\
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__2426\,
            I => \N__2423\
        );

    \I__458\ : InMux
    port map (
            O => \N__2423\,
            I => \N__2418\
        );

    \I__457\ : InMux
    port map (
            O => \N__2422\,
            I => \N__2415\
        );

    \I__456\ : InMux
    port map (
            O => \N__2421\,
            I => \N__2412\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__2418\,
            I => \Debounce_Sw1.r_CountZ0Z_6\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2415\,
            I => \Debounce_Sw1.r_CountZ0Z_6\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__2412\,
            I => \Debounce_Sw1.r_CountZ0Z_6\
        );

    \I__452\ : InMux
    port map (
            O => \N__2405\,
            I => \N__2402\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__2402\,
            I => \N__2398\
        );

    \I__450\ : InMux
    port map (
            O => \N__2401\,
            I => \N__2395\
        );

    \I__449\ : Odrv4
    port map (
            O => \N__2398\,
            I => \Debounce_Sw1.un9_r_count_9\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__2395\,
            I => \Debounce_Sw1.un9_r_count_9\
        );

    \I__447\ : InMux
    port map (
            O => \N__2390\,
            I => \N__2385\
        );

    \I__446\ : InMux
    port map (
            O => \N__2389\,
            I => \N__2382\
        );

    \I__445\ : InMux
    port map (
            O => \N__2388\,
            I => \N__2379\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2385\,
            I => \Debounce_Sw1.r_CountZ0Z_12\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2382\,
            I => \Debounce_Sw1.r_CountZ0Z_12\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__2379\,
            I => \Debounce_Sw1.r_CountZ0Z_12\
        );

    \I__441\ : InMux
    port map (
            O => \N__2372\,
            I => \N__2367\
        );

    \I__440\ : InMux
    port map (
            O => \N__2371\,
            I => \N__2364\
        );

    \I__439\ : InMux
    port map (
            O => \N__2370\,
            I => \N__2361\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2367\,
            I => \Debounce_Sw1.r_CountZ0Z_14\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__2364\,
            I => \Debounce_Sw1.r_CountZ0Z_14\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2361\,
            I => \Debounce_Sw1.r_CountZ0Z_14\
        );

    \I__435\ : CascadeMux
    port map (
            O => \N__2354\,
            I => \N__2350\
        );

    \I__434\ : InMux
    port map (
            O => \N__2353\,
            I => \N__2346\
        );

    \I__433\ : InMux
    port map (
            O => \N__2350\,
            I => \N__2343\
        );

    \I__432\ : InMux
    port map (
            O => \N__2349\,
            I => \N__2340\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2346\,
            I => \Debounce_Sw1.r_CountZ0Z_15\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2343\,
            I => \Debounce_Sw1.r_CountZ0Z_15\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2340\,
            I => \Debounce_Sw1.r_CountZ0Z_15\
        );

    \I__428\ : InMux
    port map (
            O => \N__2333\,
            I => \N__2328\
        );

    \I__427\ : InMux
    port map (
            O => \N__2332\,
            I => \N__2325\
        );

    \I__426\ : InMux
    port map (
            O => \N__2331\,
            I => \N__2322\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2328\,
            I => \Debounce_Sw1.r_CountZ0Z_7\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__2325\,
            I => \Debounce_Sw1.r_CountZ0Z_7\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2322\,
            I => \Debounce_Sw1.r_CountZ0Z_7\
        );

    \I__422\ : InMux
    port map (
            O => \N__2315\,
            I => \N__2312\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2312\,
            I => \N__2309\
        );

    \I__420\ : Odrv12
    port map (
            O => \N__2309\,
            I => \Debounce_Sw1.un9_r_count_10\
        );

    \I__419\ : InMux
    port map (
            O => \N__2306\,
            I => \N__2301\
        );

    \I__418\ : InMux
    port map (
            O => \N__2305\,
            I => \N__2298\
        );

    \I__417\ : InMux
    port map (
            O => \N__2304\,
            I => \N__2295\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2301\,
            I => \Debounce_Sw1.r_CountZ0Z_9\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2298\,
            I => \Debounce_Sw1.r_CountZ0Z_9\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2295\,
            I => \Debounce_Sw1.r_CountZ0Z_9\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__2288\,
            I => \Debounce_Sw1.un9_r_count_5_cascade_\
        );

    \I__412\ : InMux
    port map (
            O => \N__2285\,
            I => \N__2280\
        );

    \I__411\ : InMux
    port map (
            O => \N__2284\,
            I => \N__2277\
        );

    \I__410\ : InMux
    port map (
            O => \N__2283\,
            I => \N__2274\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2280\,
            I => \Debounce_Sw1.r_CountZ0Z_10\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2277\,
            I => \Debounce_Sw1.r_CountZ0Z_10\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2274\,
            I => \Debounce_Sw1.r_CountZ0Z_10\
        );

    \I__406\ : InMux
    port map (
            O => \N__2267\,
            I => \N__2264\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2264\,
            I => \Debounce_Sw1.un9_r_count_9_0\
        );

    \I__404\ : InMux
    port map (
            O => \N__2261\,
            I => \N__2258\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2258\,
            I => \N__2255\
        );

    \I__402\ : Span4Mux_h
    port map (
            O => \N__2255\,
            I => \N__2251\
        );

    \I__401\ : InMux
    port map (
            O => \N__2254\,
            I => \N__2248\
        );

    \I__400\ : Sp12to4
    port map (
            O => \N__2251\,
            I => \N__2243\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2248\,
            I => \N__2243\
        );

    \I__398\ : Span12Mux_v
    port map (
            O => \N__2243\,
            I => \N__2240\
        );

    \I__397\ : Odrv12
    port map (
            O => \N__2240\,
            I => \i_Switch_1_c\
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__2237\,
            I => \Debounce_Sw1.un9_r_count_10_0_cascade_\
        );

    \I__395\ : InMux
    port map (
            O => \N__2234\,
            I => \N__2229\
        );

    \I__394\ : InMux
    port map (
            O => \N__2233\,
            I => \N__2226\
        );

    \I__393\ : InMux
    port map (
            O => \N__2232\,
            I => \N__2223\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2229\,
            I => \N__2220\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2226\,
            I => \Debounce_Sw1.r_CountZ0Z_16\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__2223\,
            I => \Debounce_Sw1.r_CountZ0Z_16\
        );

    \I__389\ : Odrv4
    port map (
            O => \N__2220\,
            I => \Debounce_Sw1.r_CountZ0Z_16\
        );

    \I__388\ : InMux
    port map (
            O => \N__2213\,
            I => \N__2208\
        );

    \I__387\ : InMux
    port map (
            O => \N__2212\,
            I => \N__2205\
        );

    \I__386\ : InMux
    port map (
            O => \N__2211\,
            I => \N__2202\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2208\,
            I => \Debounce_Sw1.r_CountZ0Z_13\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__2205\,
            I => \Debounce_Sw1.r_CountZ0Z_13\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2202\,
            I => \Debounce_Sw1.r_CountZ0Z_13\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__2195\,
            I => \N__2191\
        );

    \I__381\ : CascadeMux
    port map (
            O => \N__2194\,
            I => \N__2187\
        );

    \I__380\ : InMux
    port map (
            O => \N__2191\,
            I => \N__2184\
        );

    \I__379\ : InMux
    port map (
            O => \N__2190\,
            I => \N__2181\
        );

    \I__378\ : InMux
    port map (
            O => \N__2187\,
            I => \N__2178\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2184\,
            I => \N__2175\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__2181\,
            I => \Debounce_Sw1.r_CountZ0Z_17\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2178\,
            I => \Debounce_Sw1.r_CountZ0Z_17\
        );

    \I__374\ : Odrv4
    port map (
            O => \N__2175\,
            I => \Debounce_Sw1.r_CountZ0Z_17\
        );

    \I__373\ : CascadeMux
    port map (
            O => \N__2168\,
            I => \N__2163\
        );

    \I__372\ : InMux
    port map (
            O => \N__2167\,
            I => \N__2160\
        );

    \I__371\ : InMux
    port map (
            O => \N__2166\,
            I => \N__2157\
        );

    \I__370\ : InMux
    port map (
            O => \N__2163\,
            I => \N__2154\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__2160\,
            I => \Debounce_Sw1.r_CountZ0Z_11\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2157\,
            I => \Debounce_Sw1.r_CountZ0Z_11\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2154\,
            I => \Debounce_Sw1.r_CountZ0Z_11\
        );

    \I__366\ : InMux
    port map (
            O => \N__2147\,
            I => \N__2144\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2144\,
            I => \Debounce_Sw1.un9_r_count_6\
        );

    \I__364\ : InMux
    port map (
            O => \N__2141\,
            I => \N__2138\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__2138\,
            I => \N__2135\
        );

    \I__362\ : Odrv4
    port map (
            O => \N__2135\,
            I => \Count_And_Toggle.r_Counter_RNO_0Z0Z_9\
        );

    \I__361\ : CascadeMux
    port map (
            O => \N__2132\,
            I => \N__2128\
        );

    \I__360\ : InMux
    port map (
            O => \N__2131\,
            I => \N__2125\
        );

    \I__359\ : InMux
    port map (
            O => \N__2128\,
            I => \N__2122\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2125\,
            I => \N__2119\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2122\,
            I => \Count_And_Toggle.r_CounterZ0Z_9\
        );

    \I__356\ : Odrv4
    port map (
            O => \N__2119\,
            I => \Count_And_Toggle.r_CounterZ0Z_9\
        );

    \I__355\ : CascadeMux
    port map (
            O => \N__2114\,
            I => \N__2111\
        );

    \I__354\ : InMux
    port map (
            O => \N__2111\,
            I => \N__2106\
        );

    \I__353\ : CascadeMux
    port map (
            O => \N__2110\,
            I => \N__2101\
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__2109\,
            I => \N__2097\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2106\,
            I => \N__2094\
        );

    \I__350\ : InMux
    port map (
            O => \N__2105\,
            I => \N__2091\
        );

    \I__349\ : CascadeMux
    port map (
            O => \N__2104\,
            I => \N__2087\
        );

    \I__348\ : InMux
    port map (
            O => \N__2101\,
            I => \N__2078\
        );

    \I__347\ : InMux
    port map (
            O => \N__2100\,
            I => \N__2078\
        );

    \I__346\ : InMux
    port map (
            O => \N__2097\,
            I => \N__2078\
        );

    \I__345\ : Span4Mux_v
    port map (
            O => \N__2094\,
            I => \N__2073\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__2091\,
            I => \N__2073\
        );

    \I__343\ : InMux
    port map (
            O => \N__2090\,
            I => \N__2070\
        );

    \I__342\ : InMux
    port map (
            O => \N__2087\,
            I => \N__2065\
        );

    \I__341\ : InMux
    port map (
            O => \N__2086\,
            I => \N__2065\
        );

    \I__340\ : InMux
    port map (
            O => \N__2085\,
            I => \N__2062\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__2078\,
            I => \Count_And_Toggle.un4_i_enable_16\
        );

    \I__338\ : Odrv4
    port map (
            O => \N__2073\,
            I => \Count_And_Toggle.un4_i_enable_16\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2070\,
            I => \Count_And_Toggle.un4_i_enable_16\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2065\,
            I => \Count_And_Toggle.un4_i_enable_16\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__2062\,
            I => \Count_And_Toggle.un4_i_enable_16\
        );

    \I__334\ : CascadeMux
    port map (
            O => \N__2051\,
            I => \N__2045\
        );

    \I__333\ : InMux
    port map (
            O => \N__2050\,
            I => \N__2038\
        );

    \I__332\ : InMux
    port map (
            O => \N__2049\,
            I => \N__2035\
        );

    \I__331\ : InMux
    port map (
            O => \N__2048\,
            I => \N__2028\
        );

    \I__330\ : InMux
    port map (
            O => \N__2045\,
            I => \N__2028\
        );

    \I__329\ : InMux
    port map (
            O => \N__2044\,
            I => \N__2028\
        );

    \I__328\ : InMux
    port map (
            O => \N__2043\,
            I => \N__2025\
        );

    \I__327\ : InMux
    port map (
            O => \N__2042\,
            I => \N__2020\
        );

    \I__326\ : InMux
    port map (
            O => \N__2041\,
            I => \N__2020\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2038\,
            I => \Count_And_Toggle.un4_i_enable_15\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2035\,
            I => \Count_And_Toggle.un4_i_enable_15\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2028\,
            I => \Count_And_Toggle.un4_i_enable_15\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__2025\,
            I => \Count_And_Toggle.un4_i_enable_15\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__2020\,
            I => \Count_And_Toggle.un4_i_enable_15\
        );

    \I__320\ : InMux
    port map (
            O => \N__2009\,
            I => \N__2006\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2006\,
            I => \Count_And_Toggle.r_Counter_RNO_0Z0Z_11\
        );

    \I__318\ : InMux
    port map (
            O => \N__2003\,
            I => \N__1999\
        );

    \I__317\ : InMux
    port map (
            O => \N__2002\,
            I => \N__1996\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__1999\,
            I => \Count_And_Toggle.r_CounterZ0Z_3\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__1996\,
            I => \Count_And_Toggle.r_CounterZ0Z_3\
        );

    \I__314\ : InMux
    port map (
            O => \N__1991\,
            I => \N__1987\
        );

    \I__313\ : InMux
    port map (
            O => \N__1990\,
            I => \N__1984\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__1987\,
            I => \Count_And_Toggle.r_CounterZ0Z_2\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__1984\,
            I => \Count_And_Toggle.r_CounterZ0Z_2\
        );

    \I__310\ : InMux
    port map (
            O => \N__1979\,
            I => \N__1972\
        );

    \I__309\ : InMux
    port map (
            O => \N__1978\,
            I => \N__1972\
        );

    \I__308\ : InMux
    port map (
            O => \N__1977\,
            I => \N__1969\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__1972\,
            I => \Count_And_Toggle.r_CounterZ0Z_1\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__1969\,
            I => \Count_And_Toggle.r_CounterZ0Z_1\
        );

    \I__305\ : InMux
    port map (
            O => \N__1964\,
            I => \N__1961\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__1961\,
            I => \N__1958\
        );

    \I__303\ : Odrv4
    port map (
            O => \N__1958\,
            I => \Count_And_Toggle.r_Counter_RNO_0Z0Z_6\
        );

    \I__302\ : CascadeMux
    port map (
            O => \N__1955\,
            I => \N__1952\
        );

    \I__301\ : InMux
    port map (
            O => \N__1952\,
            I => \N__1948\
        );

    \I__300\ : InMux
    port map (
            O => \N__1951\,
            I => \N__1945\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__1948\,
            I => \Count_And_Toggle.r_CounterZ0Z_6\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__1945\,
            I => \Count_And_Toggle.r_CounterZ0Z_6\
        );

    \I__297\ : InMux
    port map (
            O => \N__1940\,
            I => \N__1937\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__1937\,
            I => \Count_And_Toggle.r_Counter_RNO_0Z0Z_19\
        );

    \I__295\ : CascadeMux
    port map (
            O => \N__1934\,
            I => \N__1930\
        );

    \I__294\ : CascadeMux
    port map (
            O => \N__1933\,
            I => \N__1927\
        );

    \I__293\ : InMux
    port map (
            O => \N__1930\,
            I => \N__1924\
        );

    \I__292\ : InMux
    port map (
            O => \N__1927\,
            I => \N__1921\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__1924\,
            I => \Count_And_Toggle.r_CounterZ0Z_19\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__1921\,
            I => \Count_And_Toggle.r_CounterZ0Z_19\
        );

    \I__289\ : InMux
    port map (
            O => \N__1916\,
            I => \N__1912\
        );

    \I__288\ : InMux
    port map (
            O => \N__1915\,
            I => \N__1909\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__1912\,
            I => \Count_And_Toggle.r_CounterZ0Z_11\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__1909\,
            I => \Count_And_Toggle.r_CounterZ0Z_11\
        );

    \I__285\ : CascadeMux
    port map (
            O => \N__1904\,
            I => \Count_And_Toggle.un4_i_enable_15_cascade_\
        );

    \I__284\ : InMux
    port map (
            O => \N__1901\,
            I => \N__1898\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__1898\,
            I => \Count_And_Toggle.r_Counter_RNO_0Z0Z_18\
        );

    \I__282\ : InMux
    port map (
            O => \N__1895\,
            I => \N__1891\
        );

    \I__281\ : InMux
    port map (
            O => \N__1894\,
            I => \N__1888\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__1891\,
            I => \Count_And_Toggle.r_CounterZ0Z_18\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__1888\,
            I => \Count_And_Toggle.r_CounterZ0Z_18\
        );

    \I__278\ : InMux
    port map (
            O => \N__1883\,
            I => \N__1879\
        );

    \I__277\ : InMux
    port map (
            O => \N__1882\,
            I => \N__1876\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__1879\,
            I => \Count_And_Toggle.r_CounterZ0Z_15\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__1876\,
            I => \Count_And_Toggle.r_CounterZ0Z_15\
        );

    \I__274\ : InMux
    port map (
            O => \N__1871\,
            I => \N__1867\
        );

    \I__273\ : InMux
    port map (
            O => \N__1870\,
            I => \N__1864\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__1867\,
            I => \Count_And_Toggle.r_CounterZ0Z_16\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__1864\,
            I => \Count_And_Toggle.r_CounterZ0Z_16\
        );

    \I__270\ : CascadeMux
    port map (
            O => \N__1859\,
            I => \N__1853\
        );

    \I__269\ : InMux
    port map (
            O => \N__1858\,
            I => \N__1848\
        );

    \I__268\ : InMux
    port map (
            O => \N__1857\,
            I => \N__1848\
        );

    \I__267\ : InMux
    port map (
            O => \N__1856\,
            I => \N__1845\
        );

    \I__266\ : InMux
    port map (
            O => \N__1853\,
            I => \N__1842\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__1848\,
            I => \Count_And_Toggle.r_CounterZ0Z_0\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__1845\,
            I => \Count_And_Toggle.r_CounterZ0Z_0\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__1842\,
            I => \Count_And_Toggle.r_CounterZ0Z_0\
        );

    \I__262\ : InMux
    port map (
            O => \N__1835\,
            I => \N__1832\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__1832\,
            I => \Count_And_Toggle.un4_i_enable_14\
        );

    \I__260\ : InMux
    port map (
            O => \N__1829\,
            I => \N__1826\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__1826\,
            I => \Count_And_Toggle.un4_i_enable_12\
        );

    \I__258\ : CascadeMux
    port map (
            O => \N__1823\,
            I => \Count_And_Toggle.un4_i_enable_11_cascade_\
        );

    \I__257\ : InMux
    port map (
            O => \N__1820\,
            I => \N__1817\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__1817\,
            I => \Count_And_Toggle.un4_i_enable_13\
        );

    \I__255\ : InMux
    port map (
            O => \N__1814\,
            I => \Debounce_Sw1.un2_r_count_cry_13\
        );

    \I__254\ : InMux
    port map (
            O => \N__1811\,
            I => \Debounce_Sw1.un2_r_count_cry_14\
        );

    \I__253\ : InMux
    port map (
            O => \N__1808\,
            I => \Debounce_Sw1.un2_r_count_cry_15\
        );

    \I__252\ : InMux
    port map (
            O => \N__1805\,
            I => \bfn_5_7_0_\
        );

    \I__251\ : SRMux
    port map (
            O => \N__1802\,
            I => \N__1790\
        );

    \I__250\ : SRMux
    port map (
            O => \N__1801\,
            I => \N__1790\
        );

    \I__249\ : SRMux
    port map (
            O => \N__1800\,
            I => \N__1790\
        );

    \I__248\ : SRMux
    port map (
            O => \N__1799\,
            I => \N__1790\
        );

    \I__247\ : GlobalMux
    port map (
            O => \N__1790\,
            I => \N__1787\
        );

    \I__246\ : gio2CtrlBuf
    port map (
            O => \N__1787\,
            I => \Debounce_Sw1.r_count15_i_g\
        );

    \I__245\ : InMux
    port map (
            O => \N__1784\,
            I => \N__1781\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__1781\,
            I => \N__1777\
        );

    \I__243\ : InMux
    port map (
            O => \N__1780\,
            I => \N__1774\
        );

    \I__242\ : Odrv4
    port map (
            O => \N__1777\,
            I => \Count_And_Toggle.r_CounterZ0Z_12\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__1774\,
            I => \Count_And_Toggle.r_CounterZ0Z_12\
        );

    \I__240\ : InMux
    port map (
            O => \N__1769\,
            I => \N__1765\
        );

    \I__239\ : InMux
    port map (
            O => \N__1768\,
            I => \N__1762\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__1765\,
            I => \Count_And_Toggle.r_CounterZ0Z_10\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__1762\,
            I => \Count_And_Toggle.r_CounterZ0Z_10\
        );

    \I__236\ : CascadeMux
    port map (
            O => \N__1757\,
            I => \N__1754\
        );

    \I__235\ : InMux
    port map (
            O => \N__1754\,
            I => \N__1750\
        );

    \I__234\ : InMux
    port map (
            O => \N__1753\,
            I => \N__1747\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__1750\,
            I => \Count_And_Toggle.r_CounterZ0Z_13\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__1747\,
            I => \Count_And_Toggle.r_CounterZ0Z_13\
        );

    \I__231\ : InMux
    port map (
            O => \N__1742\,
            I => \N__1738\
        );

    \I__230\ : InMux
    port map (
            O => \N__1741\,
            I => \N__1735\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__1738\,
            I => \Count_And_Toggle.r_CounterZ0Z_7\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__1735\,
            I => \Count_And_Toggle.r_CounterZ0Z_7\
        );

    \I__227\ : InMux
    port map (
            O => \N__1730\,
            I => \N__1727\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1727\,
            I => \Count_And_Toggle.r_Counter_RNO_0Z0Z_8\
        );

    \I__225\ : CascadeMux
    port map (
            O => \N__1724\,
            I => \N__1720\
        );

    \I__224\ : InMux
    port map (
            O => \N__1723\,
            I => \N__1717\
        );

    \I__223\ : InMux
    port map (
            O => \N__1720\,
            I => \N__1714\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__1717\,
            I => \Count_And_Toggle.r_CounterZ0Z_8\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__1714\,
            I => \Count_And_Toggle.r_CounterZ0Z_8\
        );

    \I__220\ : InMux
    port map (
            O => \N__1709\,
            I => \N__1705\
        );

    \I__219\ : InMux
    port map (
            O => \N__1708\,
            I => \N__1702\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1705\,
            I => \Count_And_Toggle.r_CounterZ0Z_5\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__1702\,
            I => \Count_And_Toggle.r_CounterZ0Z_5\
        );

    \I__216\ : InMux
    port map (
            O => \N__1697\,
            I => \N__1693\
        );

    \I__215\ : InMux
    port map (
            O => \N__1696\,
            I => \N__1690\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__1693\,
            I => \Count_And_Toggle.r_CounterZ0Z_4\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__1690\,
            I => \Count_And_Toggle.r_CounterZ0Z_4\
        );

    \I__212\ : InMux
    port map (
            O => \N__1685\,
            I => \N__1681\
        );

    \I__211\ : InMux
    port map (
            O => \N__1684\,
            I => \N__1678\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__1681\,
            I => \Debounce_Sw1.r_CountZ0Z_5\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__1678\,
            I => \Debounce_Sw1.r_CountZ0Z_5\
        );

    \I__208\ : InMux
    port map (
            O => \N__1673\,
            I => \Debounce_Sw1.un2_r_count_cry_4\
        );

    \I__207\ : InMux
    port map (
            O => \N__1670\,
            I => \Debounce_Sw1.un2_r_count_cry_5\
        );

    \I__206\ : InMux
    port map (
            O => \N__1667\,
            I => \Debounce_Sw1.un2_r_count_cry_6\
        );

    \I__205\ : InMux
    port map (
            O => \N__1664\,
            I => \Debounce_Sw1.un2_r_count_cry_7\
        );

    \I__204\ : InMux
    port map (
            O => \N__1661\,
            I => \bfn_5_6_0_\
        );

    \I__203\ : InMux
    port map (
            O => \N__1658\,
            I => \Debounce_Sw1.un2_r_count_cry_9\
        );

    \I__202\ : InMux
    port map (
            O => \N__1655\,
            I => \Debounce_Sw1.un2_r_count_cry_10\
        );

    \I__201\ : InMux
    port map (
            O => \N__1652\,
            I => \Debounce_Sw1.un2_r_count_cry_11\
        );

    \I__200\ : InMux
    port map (
            O => \N__1649\,
            I => \Debounce_Sw1.un2_r_count_cry_12\
        );

    \I__199\ : InMux
    port map (
            O => \N__1646\,
            I => \Count_And_Toggle.un2_r_counter_cry_19\
        );

    \I__198\ : InMux
    port map (
            O => \N__1643\,
            I => \Count_And_Toggle.un2_r_counter_cry_20\
        );

    \I__197\ : InMux
    port map (
            O => \N__1640\,
            I => \Count_And_Toggle.un2_r_counter_cry_21\
        );

    \I__196\ : CascadeMux
    port map (
            O => \N__1637\,
            I => \Count_And_Toggle.r_Counter_RNO_0Z0Z_22_cascade_\
        );

    \I__195\ : InMux
    port map (
            O => \N__1634\,
            I => \N__1628\
        );

    \I__194\ : InMux
    port map (
            O => \N__1633\,
            I => \N__1628\
        );

    \I__193\ : LocalMux
    port map (
            O => \N__1628\,
            I => \Count_And_Toggle.r_CounterZ0Z_17\
        );

    \I__192\ : InMux
    port map (
            O => \N__1625\,
            I => \N__1619\
        );

    \I__191\ : InMux
    port map (
            O => \N__1624\,
            I => \N__1619\
        );

    \I__190\ : LocalMux
    port map (
            O => \N__1619\,
            I => \Count_And_Toggle.r_CounterZ0Z_22\
        );

    \I__189\ : CascadeMux
    port map (
            O => \N__1616\,
            I => \N__1613\
        );

    \I__188\ : InMux
    port map (
            O => \N__1613\,
            I => \N__1607\
        );

    \I__187\ : InMux
    port map (
            O => \N__1612\,
            I => \N__1607\
        );

    \I__186\ : LocalMux
    port map (
            O => \N__1607\,
            I => \Count_And_Toggle.r_CounterZ0Z_21\
        );

    \I__185\ : InMux
    port map (
            O => \N__1604\,
            I => \N__1598\
        );

    \I__184\ : InMux
    port map (
            O => \N__1603\,
            I => \N__1598\
        );

    \I__183\ : LocalMux
    port map (
            O => \N__1598\,
            I => \Count_And_Toggle.r_CounterZ0Z_20\
        );

    \I__182\ : InMux
    port map (
            O => \N__1595\,
            I => \N__1589\
        );

    \I__181\ : InMux
    port map (
            O => \N__1594\,
            I => \N__1582\
        );

    \I__180\ : InMux
    port map (
            O => \N__1593\,
            I => \N__1582\
        );

    \I__179\ : InMux
    port map (
            O => \N__1592\,
            I => \N__1582\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__1589\,
            I => \Debounce_Sw1.r_CountZ0Z_0\
        );

    \I__177\ : LocalMux
    port map (
            O => \N__1582\,
            I => \Debounce_Sw1.r_CountZ0Z_0\
        );

    \I__176\ : CascadeMux
    port map (
            O => \N__1577\,
            I => \N__1573\
        );

    \I__175\ : CascadeMux
    port map (
            O => \N__1576\,
            I => \N__1570\
        );

    \I__174\ : InMux
    port map (
            O => \N__1573\,
            I => \N__1566\
        );

    \I__173\ : InMux
    port map (
            O => \N__1570\,
            I => \N__1561\
        );

    \I__172\ : InMux
    port map (
            O => \N__1569\,
            I => \N__1561\
        );

    \I__171\ : LocalMux
    port map (
            O => \N__1566\,
            I => \Debounce_Sw1.r_CountZ0Z_1\
        );

    \I__170\ : LocalMux
    port map (
            O => \N__1561\,
            I => \Debounce_Sw1.r_CountZ0Z_1\
        );

    \I__169\ : InMux
    port map (
            O => \N__1556\,
            I => \N__1552\
        );

    \I__168\ : InMux
    port map (
            O => \N__1555\,
            I => \N__1549\
        );

    \I__167\ : LocalMux
    port map (
            O => \N__1552\,
            I => \Debounce_Sw1.r_CountZ0Z_2\
        );

    \I__166\ : LocalMux
    port map (
            O => \N__1549\,
            I => \Debounce_Sw1.r_CountZ0Z_2\
        );

    \I__165\ : InMux
    port map (
            O => \N__1544\,
            I => \Debounce_Sw1.un2_r_count_cry_1\
        );

    \I__164\ : CascadeMux
    port map (
            O => \N__1541\,
            I => \N__1537\
        );

    \I__163\ : InMux
    port map (
            O => \N__1540\,
            I => \N__1534\
        );

    \I__162\ : InMux
    port map (
            O => \N__1537\,
            I => \N__1531\
        );

    \I__161\ : LocalMux
    port map (
            O => \N__1534\,
            I => \Debounce_Sw1.r_CountZ0Z_3\
        );

    \I__160\ : LocalMux
    port map (
            O => \N__1531\,
            I => \Debounce_Sw1.r_CountZ0Z_3\
        );

    \I__159\ : InMux
    port map (
            O => \N__1526\,
            I => \Debounce_Sw1.un2_r_count_cry_2\
        );

    \I__158\ : InMux
    port map (
            O => \N__1523\,
            I => \N__1519\
        );

    \I__157\ : InMux
    port map (
            O => \N__1522\,
            I => \N__1516\
        );

    \I__156\ : LocalMux
    port map (
            O => \N__1519\,
            I => \Debounce_Sw1.r_CountZ0Z_4\
        );

    \I__155\ : LocalMux
    port map (
            O => \N__1516\,
            I => \Debounce_Sw1.r_CountZ0Z_4\
        );

    \I__154\ : InMux
    port map (
            O => \N__1511\,
            I => \Debounce_Sw1.un2_r_count_cry_3\
        );

    \I__153\ : InMux
    port map (
            O => \N__1508\,
            I => \Count_And_Toggle.un2_r_counter_cry_10\
        );

    \I__152\ : InMux
    port map (
            O => \N__1505\,
            I => \Count_And_Toggle.un2_r_counter_cry_11\
        );

    \I__151\ : InMux
    port map (
            O => \N__1502\,
            I => \Count_And_Toggle.un2_r_counter_cry_12\
        );

    \I__150\ : InMux
    port map (
            O => \N__1499\,
            I => \Count_And_Toggle.un2_r_counter_cry_13\
        );

    \I__149\ : InMux
    port map (
            O => \N__1496\,
            I => \Count_And_Toggle.un2_r_counter_cry_14\
        );

    \I__148\ : InMux
    port map (
            O => \N__1493\,
            I => \Count_And_Toggle.un2_r_counter_cry_15\
        );

    \I__147\ : InMux
    port map (
            O => \N__1490\,
            I => \bfn_4_9_0_\
        );

    \I__146\ : InMux
    port map (
            O => \N__1487\,
            I => \Count_And_Toggle.un2_r_counter_cry_17\
        );

    \I__145\ : InMux
    port map (
            O => \N__1484\,
            I => \Count_And_Toggle.un2_r_counter_cry_18\
        );

    \I__144\ : InMux
    port map (
            O => \N__1481\,
            I => \Count_And_Toggle.un2_r_counter_cry_1\
        );

    \I__143\ : InMux
    port map (
            O => \N__1478\,
            I => \Count_And_Toggle.un2_r_counter_cry_2\
        );

    \I__142\ : InMux
    port map (
            O => \N__1475\,
            I => \Count_And_Toggle.un2_r_counter_cry_3\
        );

    \I__141\ : InMux
    port map (
            O => \N__1472\,
            I => \Count_And_Toggle.un2_r_counter_cry_4\
        );

    \I__140\ : InMux
    port map (
            O => \N__1469\,
            I => \Count_And_Toggle.un2_r_counter_cry_5\
        );

    \I__139\ : InMux
    port map (
            O => \N__1466\,
            I => \Count_And_Toggle.un2_r_counter_cry_6\
        );

    \I__138\ : InMux
    port map (
            O => \N__1463\,
            I => \Count_And_Toggle.un2_r_counter_cry_7\
        );

    \I__137\ : InMux
    port map (
            O => \N__1460\,
            I => \bfn_4_8_0_\
        );

    \I__136\ : InMux
    port map (
            O => \N__1457\,
            I => \Count_And_Toggle.un2_r_counter_cry_9\
        );

    \I__135\ : CascadeMux
    port map (
            O => \N__1454\,
            I => \Debounce_Sw1.un9_r_count_10_cascade_\
        );

    \I__134\ : CascadeMux
    port map (
            O => \N__1451\,
            I => \Debounce_Sw1.un1_r_Count_1lt11_0_cascade_\
        );

    \I__133\ : InMux
    port map (
            O => \N__1448\,
            I => \N__1445\
        );

    \I__132\ : LocalMux
    port map (
            O => \N__1445\,
            I => \Debounce_Sw1.un1_r_Count_1lto11_1\
        );

    \I__131\ : CascadeMux
    port map (
            O => \N__1442\,
            I => \Debounce_Sw1.un1_r_Count_1lt17_cascade_\
        );

    \I__130\ : InMux
    port map (
            O => \N__1439\,
            I => \N__1436\
        );

    \I__129\ : LocalMux
    port map (
            O => \N__1436\,
            I => \Debounce_Sw1.un1_r_Count_1lto17_2\
        );

    \I__128\ : IoInMux
    port map (
            O => \N__1433\,
            I => \N__1430\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__1430\,
            I => \N__1427\
        );

    \I__126\ : Span4Mux_s3_h
    port map (
            O => \N__1427\,
            I => \N__1424\
        );

    \I__125\ : Odrv4
    port map (
            O => \N__1424\,
            I => \Debounce_Sw1.r_count15_i\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Debounce_Sw2.un2_r_count_cry_8\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Debounce_Sw2.un2_r_count_cry_16\,
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_5_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_5_0_\
        );

    \IN_MUX_bfv_5_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Debounce_Sw1.un2_r_count_cry_8\,
            carryinitout => \bfn_5_6_0_\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Debounce_Sw1.un2_r_count_cry_16\,
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_4_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_7_0_\
        );

    \IN_MUX_bfv_4_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Count_And_Toggle.un2_r_counter_cry_8\,
            carryinitout => \bfn_4_8_0_\
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Count_And_Toggle.un2_r_counter_cry_16\,
            carryinitout => \bfn_4_9_0_\
        );

    \Debounce_Sw2.r_State_e_0_RNIK82U4_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2495\,
            GLOBALBUFFEROUTPUT => \Debounce_Sw2.N_9_g\
        );

    \Debounce_Sw1.r_State_RNIDSE73_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1433\,
            GLOBALBUFFEROUTPUT => \Debounce_Sw1.r_count15_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \Debounce_Sw1.r_Count_RNI720A_4_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1522\,
            in2 => \_gnd_net_\,
            in3 => \N__1684\,
            lcout => \Debounce_Sw1.un9_r_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.r_Count_RNIGFOJ_10_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2283\,
            in1 => \N__2304\,
            in2 => \N__2168\,
            in3 => \N__2442\,
            lcout => \Debounce_Sw1.un1_r_Count_1lto11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.r_Count_RNIMUGJ_17_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2234\,
            in1 => \N__2349\,
            in2 => \N__2195\,
            in3 => \N__2370\,
            lcout => \Debounce_Sw1.un1_r_Count_1lto17_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.r_Count_1_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1576\,
            in3 => \N__1593\,
            lcout => \Debounce_Sw1.r_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3075\,
            ce => 'H',
            sr => \N__1799\
        );

    \Debounce_Sw1.r_Count_RNI2OVJ_1_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1592\,
            in1 => \N__1569\,
            in2 => \N__1541\,
            in3 => \N__1555\,
            lcout => \Debounce_Sw1.un9_r_count_10\,
            ltout => \Debounce_Sw1.un9_r_count_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.r_Count_RNIK0081_6_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010101010"
        )
    port map (
            in0 => \N__2331\,
            in1 => \N__2421\,
            in2 => \N__1454\,
            in3 => \N__2401\,
            lcout => OPEN,
            ltout => \Debounce_Sw1.un1_r_Count_1lt11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.r_Count_RNI9PG52_12_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100010001"
        )
    port map (
            in0 => \N__2211\,
            in1 => \N__2388\,
            in2 => \N__1451\,
            in3 => \N__1448\,
            lcout => OPEN,
            ltout => \Debounce_Sw1.un1_r_Count_1lt17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.r_State_RNIDSE73_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110011001"
        )
    port map (
            in0 => \N__2261\,
            in1 => \N__2974\,
            in2 => \N__1442\,
            in3 => \N__1439\,
            lcout => \Debounce_Sw1.r_count15_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.r_Count_0_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__1594\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Debounce_Sw1.r_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3075\,
            ce => 'H',
            sr => \N__1799\
        );

    \Count_And_Toggle.un2_r_counter_cry_1_c_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1977\,
            in2 => \N__1859\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_7_0_\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_2_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1990\,
            in2 => \_gnd_net_\,
            in3 => \N__1481\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_2\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_1\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_2\,
            clk => \N__3072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_3_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2002\,
            in2 => \_gnd_net_\,
            in3 => \N__1478\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_3\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_2\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_3\,
            clk => \N__3072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_4_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1696\,
            in2 => \_gnd_net_\,
            in3 => \N__1475\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_4\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_3\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_4\,
            clk => \N__3072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_5_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1708\,
            in2 => \_gnd_net_\,
            in3 => \N__1472\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_5\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_4\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_5\,
            clk => \N__3072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNO_0_6_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1951\,
            in2 => \_gnd_net_\,
            in3 => \N__1469\,
            lcout => \Count_And_Toggle.r_Counter_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_5\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_7_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1741\,
            in2 => \_gnd_net_\,
            in3 => \N__1466\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_7\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_6\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_7\,
            clk => \N__3072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNO_0_8_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1724\,
            in3 => \N__1463\,
            lcout => \Count_And_Toggle.r_Counter_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_7\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNO_0_9_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2131\,
            in2 => \_gnd_net_\,
            in3 => \N__1460\,
            lcout => \Count_And_Toggle.r_Counter_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_4_8_0_\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_10_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1768\,
            in2 => \_gnd_net_\,
            in3 => \N__1457\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_10\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_9\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_10\,
            clk => \N__3070\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNO_0_11_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1915\,
            in2 => \_gnd_net_\,
            in3 => \N__1508\,
            lcout => \Count_And_Toggle.r_Counter_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_10\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_12_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1780\,
            in2 => \_gnd_net_\,
            in3 => \N__1505\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_12\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_11\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_12\,
            clk => \N__3070\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_13_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1753\,
            in2 => \_gnd_net_\,
            in3 => \N__1502\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_13\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_12\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_13\,
            clk => \N__3070\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNO_0_14_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2455\,
            in2 => \_gnd_net_\,
            in3 => \N__1499\,
            lcout => \Count_And_Toggle.r_Counter_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_13\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_15_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1882\,
            in2 => \_gnd_net_\,
            in3 => \N__1496\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_15\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_14\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_15\,
            clk => \N__3070\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_16_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1870\,
            in2 => \_gnd_net_\,
            in3 => \N__1493\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_16\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_15\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_16\,
            clk => \N__3070\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_17_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1633\,
            in2 => \_gnd_net_\,
            in3 => \N__1490\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_17\,
            clk => \N__3073\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNO_0_18_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1894\,
            in2 => \_gnd_net_\,
            in3 => \N__1487\,
            lcout => \Count_And_Toggle.r_Counter_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_17\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNO_0_19_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1933\,
            in3 => \N__1484\,
            lcout => \Count_And_Toggle.r_Counter_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_18\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_20_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1603\,
            in2 => \_gnd_net_\,
            in3 => \N__1646\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_20\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_19\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_20\,
            clk => \N__3073\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_21_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1612\,
            in2 => \_gnd_net_\,
            in3 => \N__1643\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_21\,
            ltout => OPEN,
            carryin => \Count_And_Toggle.un2_r_counter_cry_20\,
            carryout => \Count_And_Toggle.un2_r_counter_cry_21\,
            clk => \N__3073\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNO_0_22_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1625\,
            in2 => \_gnd_net_\,
            in3 => \N__1640\,
            lcout => OPEN,
            ltout => \Count_And_Toggle.r_Counter_RNO_0Z0Z_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_22_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__2085\,
            in1 => \N__2049\,
            in2 => \N__1637\,
            in3 => \N__2572\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3073\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNITEQL1_22_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__1634\,
            in1 => \N__1624\,
            in2 => \N__1616\,
            in3 => \N__1604\,
            lcout => \Count_And_Toggle.un4_i_enable_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.un2_r_count_cry_1_c_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1595\,
            in2 => \N__1577\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_5_0_\,
            carryout => \Debounce_Sw1.un2_r_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.r_Count_2_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1556\,
            in2 => \_gnd_net_\,
            in3 => \N__1544\,
            lcout => \Debounce_Sw1.r_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_1\,
            carryout => \Debounce_Sw1.un2_r_count_cry_2\,
            clk => \N__3081\,
            ce => 'H',
            sr => \N__1802\
        );

    \Debounce_Sw1.r_Count_3_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1540\,
            in2 => \_gnd_net_\,
            in3 => \N__1526\,
            lcout => \Debounce_Sw1.r_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_2\,
            carryout => \Debounce_Sw1.un2_r_count_cry_3\,
            clk => \N__3081\,
            ce => 'H',
            sr => \N__1802\
        );

    \Debounce_Sw1.r_Count_4_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1523\,
            in2 => \_gnd_net_\,
            in3 => \N__1511\,
            lcout => \Debounce_Sw1.r_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_3\,
            carryout => \Debounce_Sw1.un2_r_count_cry_4\,
            clk => \N__3081\,
            ce => 'H',
            sr => \N__1802\
        );

    \Debounce_Sw1.r_Count_5_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1685\,
            in2 => \_gnd_net_\,
            in3 => \N__1673\,
            lcout => \Debounce_Sw1.r_CountZ0Z_5\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_4\,
            carryout => \Debounce_Sw1.un2_r_count_cry_5\,
            clk => \N__3081\,
            ce => 'H',
            sr => \N__1802\
        );

    \Debounce_Sw1.r_Count_6_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2422\,
            in2 => \_gnd_net_\,
            in3 => \N__1670\,
            lcout => \Debounce_Sw1.r_CountZ0Z_6\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_5\,
            carryout => \Debounce_Sw1.un2_r_count_cry_6\,
            clk => \N__3081\,
            ce => 'H',
            sr => \N__1802\
        );

    \Debounce_Sw1.r_Count_7_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2333\,
            in2 => \_gnd_net_\,
            in3 => \N__1667\,
            lcout => \Debounce_Sw1.r_CountZ0Z_7\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_6\,
            carryout => \Debounce_Sw1.un2_r_count_cry_7\,
            clk => \N__3081\,
            ce => 'H',
            sr => \N__1802\
        );

    \Debounce_Sw1.r_Count_8_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2443\,
            in2 => \_gnd_net_\,
            in3 => \N__1664\,
            lcout => \Debounce_Sw1.r_CountZ0Z_8\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_7\,
            carryout => \Debounce_Sw1.un2_r_count_cry_8\,
            clk => \N__3081\,
            ce => 'H',
            sr => \N__1802\
        );

    \Debounce_Sw1.r_Count_9_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2305\,
            in2 => \_gnd_net_\,
            in3 => \N__1661\,
            lcout => \Debounce_Sw1.r_CountZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_5_6_0_\,
            carryout => \Debounce_Sw1.un2_r_count_cry_9\,
            clk => \N__3079\,
            ce => 'H',
            sr => \N__1801\
        );

    \Debounce_Sw1.r_Count_10_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2284\,
            in2 => \_gnd_net_\,
            in3 => \N__1658\,
            lcout => \Debounce_Sw1.r_CountZ0Z_10\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_9\,
            carryout => \Debounce_Sw1.un2_r_count_cry_10\,
            clk => \N__3079\,
            ce => 'H',
            sr => \N__1801\
        );

    \Debounce_Sw1.r_Count_11_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2167\,
            in2 => \_gnd_net_\,
            in3 => \N__1655\,
            lcout => \Debounce_Sw1.r_CountZ0Z_11\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_10\,
            carryout => \Debounce_Sw1.un2_r_count_cry_11\,
            clk => \N__3079\,
            ce => 'H',
            sr => \N__1801\
        );

    \Debounce_Sw1.r_Count_12_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2390\,
            in2 => \_gnd_net_\,
            in3 => \N__1652\,
            lcout => \Debounce_Sw1.r_CountZ0Z_12\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_11\,
            carryout => \Debounce_Sw1.un2_r_count_cry_12\,
            clk => \N__3079\,
            ce => 'H',
            sr => \N__1801\
        );

    \Debounce_Sw1.r_Count_13_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2213\,
            in2 => \_gnd_net_\,
            in3 => \N__1649\,
            lcout => \Debounce_Sw1.r_CountZ0Z_13\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_12\,
            carryout => \Debounce_Sw1.un2_r_count_cry_13\,
            clk => \N__3079\,
            ce => 'H',
            sr => \N__1801\
        );

    \Debounce_Sw1.r_Count_14_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2372\,
            in2 => \_gnd_net_\,
            in3 => \N__1814\,
            lcout => \Debounce_Sw1.r_CountZ0Z_14\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_13\,
            carryout => \Debounce_Sw1.un2_r_count_cry_14\,
            clk => \N__3079\,
            ce => 'H',
            sr => \N__1801\
        );

    \Debounce_Sw1.r_Count_15_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2353\,
            in2 => \_gnd_net_\,
            in3 => \N__1811\,
            lcout => \Debounce_Sw1.r_CountZ0Z_15\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_14\,
            carryout => \Debounce_Sw1.un2_r_count_cry_15\,
            clk => \N__3079\,
            ce => 'H',
            sr => \N__1801\
        );

    \Debounce_Sw1.r_Count_16_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2233\,
            in2 => \_gnd_net_\,
            in3 => \N__1808\,
            lcout => \Debounce_Sw1.r_CountZ0Z_16\,
            ltout => OPEN,
            carryin => \Debounce_Sw1.un2_r_count_cry_15\,
            carryout => \Debounce_Sw1.un2_r_count_cry_16\,
            clk => \N__3079\,
            ce => 'H',
            sr => \N__1801\
        );

    \Debounce_Sw1.r_Count_17_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2190\,
            in2 => \_gnd_net_\,
            in3 => \N__1805\,
            lcout => \Debounce_Sw1.r_CountZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3076\,
            ce => 'H',
            sr => \N__1800\
        );

    \Count_And_Toggle.r_Counter_RNIBHPL1_10_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1784\,
            in1 => \N__1769\,
            in2 => \N__1757\,
            in3 => \N__1742\,
            lcout => \Count_And_Toggle.un4_i_enable_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_8_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2048\,
            in1 => \N__2571\,
            in2 => \N__2110\,
            in3 => \N__1730\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_1_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__1858\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1979\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_0_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1857\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNI6J0M1_4_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1723\,
            in1 => \N__1709\,
            in2 => \N__2132\,
            in3 => \N__1697\,
            lcout => \Count_And_Toggle.un4_i_enable_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_11_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2044\,
            in1 => \N__2569\,
            in2 => \N__2109\,
            in3 => \N__2009\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNIO40M1_1_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__2003\,
            in1 => \N__1991\,
            in2 => \N__1955\,
            in3 => \N__1978\,
            lcout => \Count_And_Toggle.un4_i_enable_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_6_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__2100\,
            in1 => \N__1964\,
            in2 => \N__2051\,
            in3 => \N__2570\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_19_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2567\,
            in1 => \N__2042\,
            in2 => \N__2104\,
            in3 => \N__1940\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNI6LNL1_11_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1895\,
            in1 => \N__2456\,
            in2 => \N__1934\,
            in3 => \N__1916\,
            lcout => \Count_And_Toggle.un4_i_enable_15\,
            ltout => \Count_And_Toggle.un4_i_enable_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_18_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2090\,
            in1 => \N__2566\,
            in2 => \N__1904\,
            in3 => \N__1901\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNIMOB81_15_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__1883\,
            in1 => \N__1871\,
            in2 => \_gnd_net_\,
            in3 => \N__1856\,
            lcout => OPEN,
            ltout => \Count_And_Toggle.un4_i_enable_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_RNIV16A6_10_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1835\,
            in1 => \N__1829\,
            in2 => \N__1823\,
            in3 => \N__1820\,
            lcout => \Count_And_Toggle.un4_i_enable_20\,
            ltout => \Count_And_Toggle.un4_i_enable_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_14_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2086\,
            in1 => \N__2041\,
            in2 => \N__2465\,
            in3 => \N__2462\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.r_State_RNO_0_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__2444\,
            in1 => \N__2147\,
            in2 => \N__2426\,
            in3 => \N__2405\,
            lcout => \Debounce_Sw1.un9_r_count_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.r_State_RNO_3_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2389\,
            in1 => \N__2371\,
            in2 => \N__2354\,
            in3 => \N__2332\,
            lcout => OPEN,
            ltout => \Debounce_Sw1.un9_r_count_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.r_State_RNO_1_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__2315\,
            in1 => \N__2306\,
            in2 => \N__2288\,
            in3 => \N__2285\,
            lcout => OPEN,
            ltout => \Debounce_Sw1.un9_r_count_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.r_State_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__2267\,
            in1 => \N__2254\,
            in2 => \N__2237\,
            in3 => \N__2973\,
            lcout => \w_Switch_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw1.r_State_RNO_2_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__2232\,
            in1 => \N__2212\,
            in2 => \N__2194\,
            in3 => \N__2166\,
            lcout => \Debounce_Sw1.un9_r_count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.r_Counter_9_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2050\,
            in1 => \N__2573\,
            in2 => \N__2114\,
            in3 => \N__2141\,
            lcout => \Count_And_Toggle.r_CounterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3074\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Count_And_Toggle.o_Toggle_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__2105\,
            in1 => \N__2043\,
            in2 => \N__2935\,
            in3 => \N__2568\,
            lcout => \w_Toggle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw2.r_State_e_0_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2524\,
            lcout => \w_Switch_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3082\,
            ce => \N__2474\,
            sr => \_gnd_net_\
        );

    \Debounce_Sw2.r_Count_1_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__2684\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2662\,
            lcout => \Debounce_Sw2.r_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3078\,
            ce => 'H',
            sr => \N__3028\
        );

    \Debounce_Sw2.r_Count_0_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2683\,
            lcout => \Debounce_Sw2.r_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3078\,
            ce => 'H',
            sr => \N__3028\
        );

    \Debounce_Sw2.r_Count_RNIV5631_4_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__2591\,
            in1 => \N__2605\,
            in2 => \_gnd_net_\,
            in3 => \N__2875\,
            lcout => \Debounce_Sw2.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw2.r_Count_RNI64TE1_1_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2620\,
            in1 => \N__2658\,
            in2 => \N__2642\,
            in3 => \N__2681\,
            lcout => \Debounce_Sw2.un9_r_count_10\,
            ltout => \Debounce_Sw2.un9_r_count_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw2.r_Count_RNISOQT2_7_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2856\,
            in2 => \N__2534\,
            in3 => \N__2719\,
            lcout => OPEN,
            ltout => \Debounce_Sw2.N_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw2.r_Count_RNINN314_12_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__2772\,
            in1 => \N__2754\,
            in2 => \N__2531\,
            in3 => \N__2692\,
            lcout => OPEN,
            ltout => \Debounce_Sw2.N_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw2.r_State_e_0_RNIK82U4_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011010101"
        )
    port map (
            in0 => \N__2528\,
            in1 => \N__2701\,
            in2 => \N__2498\,
            in3 => \N__2893\,
            lcout => \Debounce_Sw2.N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw2.r_State_e_0_RNO_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__2702\,
            in1 => \N__2708\,
            in2 => \N__2483\,
            in3 => \N__2693\,
            lcout => \Debounce_Sw2.r_State_e_0_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw2.r_State_e_0_RNO_0_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__2720\,
            in1 => \N__2773\,
            in2 => \N__2861\,
            in3 => \N__2755\,
            lcout => \Debounce_Sw2.un9_r_count_0_a3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw2.r_Count_RNIQEQB_17_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3121\,
            in1 => \N__3136\,
            in2 => \N__3104\,
            in3 => \N__2734\,
            lcout => \Debounce_Sw2.N_22_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw2.r_Count_RNIKTBT_10_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2806\,
            in1 => \N__2821\,
            in2 => \N__2792\,
            in3 => \N__2836\,
            lcout => \Debounce_Sw2.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw2.un2_r_count_cry_1_c_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2682\,
            in2 => \N__2663\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \Debounce_Sw2.un2_r_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Debounce_Sw2.r_Count_2_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2638\,
            in2 => \_gnd_net_\,
            in3 => \N__2624\,
            lcout => \Debounce_Sw2.r_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_1\,
            carryout => \Debounce_Sw2.un2_r_count_cry_2\,
            clk => \N__3084\,
            ce => 'H',
            sr => \N__3029\
        );

    \Debounce_Sw2.r_Count_3_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2621\,
            in2 => \_gnd_net_\,
            in3 => \N__2609\,
            lcout => \Debounce_Sw2.r_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_2\,
            carryout => \Debounce_Sw2.un2_r_count_cry_3\,
            clk => \N__3084\,
            ce => 'H',
            sr => \N__3029\
        );

    \Debounce_Sw2.r_Count_4_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2606\,
            in2 => \_gnd_net_\,
            in3 => \N__2594\,
            lcout => \Debounce_Sw2.r_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_3\,
            carryout => \Debounce_Sw2.un2_r_count_cry_4\,
            clk => \N__3084\,
            ce => 'H',
            sr => \N__3029\
        );

    \Debounce_Sw2.r_Count_5_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2590\,
            in2 => \_gnd_net_\,
            in3 => \N__2576\,
            lcout => \Debounce_Sw2.r_CountZ0Z_5\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_4\,
            carryout => \Debounce_Sw2.un2_r_count_cry_5\,
            clk => \N__3084\,
            ce => 'H',
            sr => \N__3029\
        );

    \Debounce_Sw2.r_Count_6_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2876\,
            in2 => \_gnd_net_\,
            in3 => \N__2864\,
            lcout => \Debounce_Sw2.r_CountZ0Z_6\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_5\,
            carryout => \Debounce_Sw2.un2_r_count_cry_6\,
            clk => \N__3084\,
            ce => 'H',
            sr => \N__3029\
        );

    \Debounce_Sw2.r_Count_7_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2860\,
            in2 => \_gnd_net_\,
            in3 => \N__2840\,
            lcout => \Debounce_Sw2.r_CountZ0Z_7\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_6\,
            carryout => \Debounce_Sw2.un2_r_count_cry_7\,
            clk => \N__3084\,
            ce => 'H',
            sr => \N__3029\
        );

    \Debounce_Sw2.r_Count_8_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2837\,
            in2 => \_gnd_net_\,
            in3 => \N__2825\,
            lcout => \Debounce_Sw2.r_CountZ0Z_8\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_7\,
            carryout => \Debounce_Sw2.un2_r_count_cry_8\,
            clk => \N__3084\,
            ce => 'H',
            sr => \N__3029\
        );

    \Debounce_Sw2.r_Count_9_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2822\,
            in2 => \_gnd_net_\,
            in3 => \N__2810\,
            lcout => \Debounce_Sw2.r_CountZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \Debounce_Sw2.un2_r_count_cry_9\,
            clk => \N__3085\,
            ce => 'H',
            sr => \N__3027\
        );

    \Debounce_Sw2.r_Count_10_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2807\,
            in2 => \_gnd_net_\,
            in3 => \N__2795\,
            lcout => \Debounce_Sw2.r_CountZ0Z_10\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_9\,
            carryout => \Debounce_Sw2.un2_r_count_cry_10\,
            clk => \N__3085\,
            ce => 'H',
            sr => \N__3027\
        );

    \Debounce_Sw2.r_Count_11_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2791\,
            in2 => \_gnd_net_\,
            in3 => \N__2777\,
            lcout => \Debounce_Sw2.r_CountZ0Z_11\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_10\,
            carryout => \Debounce_Sw2.un2_r_count_cry_11\,
            clk => \N__3085\,
            ce => 'H',
            sr => \N__3027\
        );

    \Debounce_Sw2.r_Count_12_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2774\,
            in2 => \_gnd_net_\,
            in3 => \N__2759\,
            lcout => \Debounce_Sw2.r_CountZ0Z_12\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_11\,
            carryout => \Debounce_Sw2.un2_r_count_cry_12\,
            clk => \N__3085\,
            ce => 'H',
            sr => \N__3027\
        );

    \Debounce_Sw2.r_Count_13_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2756\,
            in2 => \_gnd_net_\,
            in3 => \N__2738\,
            lcout => \Debounce_Sw2.r_CountZ0Z_13\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_12\,
            carryout => \Debounce_Sw2.un2_r_count_cry_13\,
            clk => \N__3085\,
            ce => 'H',
            sr => \N__3027\
        );

    \Debounce_Sw2.r_Count_14_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2735\,
            in2 => \_gnd_net_\,
            in3 => \N__2723\,
            lcout => \Debounce_Sw2.r_CountZ0Z_14\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_13\,
            carryout => \Debounce_Sw2.un2_r_count_cry_14\,
            clk => \N__3085\,
            ce => 'H',
            sr => \N__3027\
        );

    \Debounce_Sw2.r_Count_15_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3137\,
            in2 => \_gnd_net_\,
            in3 => \N__3125\,
            lcout => \Debounce_Sw2.r_CountZ0Z_15\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_14\,
            carryout => \Debounce_Sw2.un2_r_count_cry_15\,
            clk => \N__3085\,
            ce => 'H',
            sr => \N__3027\
        );

    \Debounce_Sw2.r_Count_16_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3122\,
            in2 => \_gnd_net_\,
            in3 => \N__3110\,
            lcout => \Debounce_Sw2.r_CountZ0Z_16\,
            ltout => OPEN,
            carryin => \Debounce_Sw2.un2_r_count_cry_15\,
            carryout => \Debounce_Sw2.un2_r_count_cry_16\,
            clk => \N__3085\,
            ce => 'H',
            sr => \N__3027\
        );

    \Debounce_Sw2.r_Count_17_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3100\,
            in2 => \_gnd_net_\,
            in3 => \N__3107\,
            lcout => \Debounce_Sw2.r_CountZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3086\,
            ce => 'H',
            sr => \N__3026\
        );

    \Demux.o_Data2_0_a3_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__2953\,
            in1 => \_gnd_net_\,
            in2 => \N__2918\,
            in3 => \N__2991\,
            lcout => \o_LED_2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Demux.o_Data3_0_a3_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__2992\,
            in1 => \N__2954\,
            in2 => \_gnd_net_\,
            in3 => \N__2917\,
            lcout => \o_LED_3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Demux.o_Data1_0_a3_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__2990\,
            in1 => \N__2952\,
            in2 => \_gnd_net_\,
            in3 => \N__2913\,
            lcout => \o_LED_1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Demux.o_Data4_0_a3_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2993\,
            in1 => \N__2951\,
            in2 => \_gnd_net_\,
            in3 => \N__2912\,
            lcout => \o_LED_4_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
