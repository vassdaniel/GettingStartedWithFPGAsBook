// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 20 2024 18:30:00

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Demux_Toggle_TOP" view "INTERFACE"

module Demux_Toggle_TOP (
    o_LED_3,
    o_LED_1,
    i_Switch_2,
    i_Clk,
    o_LED_4,
    o_LED_2,
    i_Switch_1);

    output o_LED_3;
    output o_LED_1;
    input i_Switch_2;
    input i_Clk;
    output o_LED_4;
    output o_LED_2;
    input i_Switch_1;

    wire N__3212;
    wire N__3211;
    wire N__3210;
    wire N__3201;
    wire N__3200;
    wire N__3199;
    wire N__3192;
    wire N__3191;
    wire N__3190;
    wire N__3183;
    wire N__3182;
    wire N__3181;
    wire N__3174;
    wire N__3173;
    wire N__3172;
    wire N__3165;
    wire N__3164;
    wire N__3163;
    wire N__3156;
    wire N__3155;
    wire N__3154;
    wire N__3137;
    wire N__3136;
    wire N__3133;
    wire N__3130;
    wire N__3125;
    wire N__3122;
    wire N__3121;
    wire N__3118;
    wire N__3115;
    wire N__3110;
    wire N__3107;
    wire N__3104;
    wire N__3101;
    wire N__3100;
    wire N__3097;
    wire N__3094;
    wire N__3091;
    wire N__3086;
    wire N__3085;
    wire N__3084;
    wire N__3083;
    wire N__3082;
    wire N__3081;
    wire N__3080;
    wire N__3079;
    wire N__3078;
    wire N__3077;
    wire N__3076;
    wire N__3075;
    wire N__3074;
    wire N__3073;
    wire N__3072;
    wire N__3071;
    wire N__3070;
    wire N__3035;
    wire N__3032;
    wire N__3029;
    wire N__3028;
    wire N__3027;
    wire N__3026;
    wire N__3017;
    wire N__3014;
    wire N__3011;
    wire N__3008;
    wire N__3005;
    wire N__3002;
    wire N__2999;
    wire N__2996;
    wire N__2993;
    wire N__2992;
    wire N__2991;
    wire N__2990;
    wire N__2987;
    wire N__2980;
    wire N__2975;
    wire N__2974;
    wire N__2973;
    wire N__2970;
    wire N__2967;
    wire N__2964;
    wire N__2959;
    wire N__2954;
    wire N__2953;
    wire N__2952;
    wire N__2951;
    wire N__2944;
    wire N__2941;
    wire N__2936;
    wire N__2935;
    wire N__2932;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2918;
    wire N__2917;
    wire N__2914;
    wire N__2913;
    wire N__2912;
    wire N__2905;
    wire N__2902;
    wire N__2897;
    wire N__2894;
    wire N__2893;
    wire N__2890;
    wire N__2887;
    wire N__2882;
    wire N__2879;
    wire N__2876;
    wire N__2875;
    wire N__2872;
    wire N__2869;
    wire N__2864;
    wire N__2861;
    wire N__2860;
    wire N__2857;
    wire N__2856;
    wire N__2853;
    wire N__2850;
    wire N__2847;
    wire N__2840;
    wire N__2837;
    wire N__2836;
    wire N__2833;
    wire N__2830;
    wire N__2825;
    wire N__2822;
    wire N__2821;
    wire N__2818;
    wire N__2815;
    wire N__2810;
    wire N__2807;
    wire N__2806;
    wire N__2803;
    wire N__2800;
    wire N__2795;
    wire N__2792;
    wire N__2791;
    wire N__2788;
    wire N__2785;
    wire N__2782;
    wire N__2777;
    wire N__2774;
    wire N__2773;
    wire N__2772;
    wire N__2769;
    wire N__2764;
    wire N__2759;
    wire N__2756;
    wire N__2755;
    wire N__2754;
    wire N__2751;
    wire N__2748;
    wire N__2745;
    wire N__2738;
    wire N__2735;
    wire N__2734;
    wire N__2731;
    wire N__2728;
    wire N__2723;
    wire N__2720;
    wire N__2719;
    wire N__2716;
    wire N__2713;
    wire N__2708;
    wire N__2705;
    wire N__2702;
    wire N__2701;
    wire N__2696;
    wire N__2693;
    wire N__2692;
    wire N__2687;
    wire N__2684;
    wire N__2683;
    wire N__2682;
    wire N__2681;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2663;
    wire N__2662;
    wire N__2659;
    wire N__2658;
    wire N__2655;
    wire N__2652;
    wire N__2649;
    wire N__2642;
    wire N__2639;
    wire N__2638;
    wire N__2635;
    wire N__2632;
    wire N__2629;
    wire N__2624;
    wire N__2621;
    wire N__2620;
    wire N__2617;
    wire N__2614;
    wire N__2609;
    wire N__2606;
    wire N__2605;
    wire N__2602;
    wire N__2599;
    wire N__2594;
    wire N__2591;
    wire N__2590;
    wire N__2587;
    wire N__2584;
    wire N__2581;
    wire N__2576;
    wire N__2573;
    wire N__2572;
    wire N__2571;
    wire N__2570;
    wire N__2569;
    wire N__2568;
    wire N__2567;
    wire N__2566;
    wire N__2563;
    wire N__2560;
    wire N__2553;
    wire N__2550;
    wire N__2545;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2525;
    wire N__2524;
    wire N__2521;
    wire N__2518;
    wire N__2515;
    wire N__2512;
    wire N__2509;
    wire N__2506;
    wire N__2503;
    wire N__2498;
    wire N__2495;
    wire N__2492;
    wire N__2489;
    wire N__2486;
    wire N__2483;
    wire N__2480;
    wire N__2477;
    wire N__2474;
    wire N__2471;
    wire N__2468;
    wire N__2465;
    wire N__2462;
    wire N__2459;
    wire N__2456;
    wire N__2455;
    wire N__2452;
    wire N__2449;
    wire N__2444;
    wire N__2443;
    wire N__2442;
    wire N__2439;
    wire N__2436;
    wire N__2433;
    wire N__2426;
    wire N__2423;
    wire N__2422;
    wire N__2421;
    wire N__2418;
    wire N__2415;
    wire N__2412;
    wire N__2405;
    wire N__2402;
    wire N__2401;
    wire N__2398;
    wire N__2395;
    wire N__2390;
    wire N__2389;
    wire N__2388;
    wire N__2385;
    wire N__2382;
    wire N__2379;
    wire N__2372;
    wire N__2371;
    wire N__2370;
    wire N__2367;
    wire N__2364;
    wire N__2361;
    wire N__2354;
    wire N__2353;
    wire N__2350;
    wire N__2349;
    wire N__2346;
    wire N__2343;
    wire N__2340;
    wire N__2333;
    wire N__2332;
    wire N__2331;
    wire N__2328;
    wire N__2325;
    wire N__2322;
    wire N__2315;
    wire N__2312;
    wire N__2309;
    wire N__2306;
    wire N__2305;
    wire N__2304;
    wire N__2301;
    wire N__2298;
    wire N__2295;
    wire N__2288;
    wire N__2285;
    wire N__2284;
    wire N__2283;
    wire N__2280;
    wire N__2277;
    wire N__2274;
    wire N__2267;
    wire N__2264;
    wire N__2261;
    wire N__2258;
    wire N__2255;
    wire N__2254;
    wire N__2251;
    wire N__2248;
    wire N__2243;
    wire N__2240;
    wire N__2237;
    wire N__2234;
    wire N__2233;
    wire N__2232;
    wire N__2229;
    wire N__2226;
    wire N__2223;
    wire N__2220;
    wire N__2213;
    wire N__2212;
    wire N__2211;
    wire N__2208;
    wire N__2205;
    wire N__2202;
    wire N__2195;
    wire N__2194;
    wire N__2191;
    wire N__2190;
    wire N__2187;
    wire N__2184;
    wire N__2181;
    wire N__2178;
    wire N__2175;
    wire N__2168;
    wire N__2167;
    wire N__2166;
    wire N__2163;
    wire N__2160;
    wire N__2157;
    wire N__2154;
    wire N__2147;
    wire N__2144;
    wire N__2141;
    wire N__2138;
    wire N__2135;
    wire N__2132;
    wire N__2131;
    wire N__2128;
    wire N__2125;
    wire N__2122;
    wire N__2119;
    wire N__2114;
    wire N__2111;
    wire N__2110;
    wire N__2109;
    wire N__2106;
    wire N__2105;
    wire N__2104;
    wire N__2101;
    wire N__2100;
    wire N__2097;
    wire N__2094;
    wire N__2091;
    wire N__2090;
    wire N__2087;
    wire N__2086;
    wire N__2085;
    wire N__2078;
    wire N__2073;
    wire N__2070;
    wire N__2065;
    wire N__2062;
    wire N__2051;
    wire N__2050;
    wire N__2049;
    wire N__2048;
    wire N__2045;
    wire N__2044;
    wire N__2043;
    wire N__2042;
    wire N__2041;
    wire N__2038;
    wire N__2035;
    wire N__2028;
    wire N__2025;
    wire N__2020;
    wire N__2009;
    wire N__2006;
    wire N__2003;
    wire N__2002;
    wire N__1999;
    wire N__1996;
    wire N__1991;
    wire N__1990;
    wire N__1987;
    wire N__1984;
    wire N__1979;
    wire N__1978;
    wire N__1977;
    wire N__1972;
    wire N__1969;
    wire N__1964;
    wire N__1961;
    wire N__1958;
    wire N__1955;
    wire N__1952;
    wire N__1951;
    wire N__1948;
    wire N__1945;
    wire N__1940;
    wire N__1937;
    wire N__1934;
    wire N__1933;
    wire N__1930;
    wire N__1927;
    wire N__1924;
    wire N__1921;
    wire N__1916;
    wire N__1915;
    wire N__1912;
    wire N__1909;
    wire N__1904;
    wire N__1901;
    wire N__1898;
    wire N__1895;
    wire N__1894;
    wire N__1891;
    wire N__1888;
    wire N__1883;
    wire N__1882;
    wire N__1879;
    wire N__1876;
    wire N__1871;
    wire N__1870;
    wire N__1867;
    wire N__1864;
    wire N__1859;
    wire N__1858;
    wire N__1857;
    wire N__1856;
    wire N__1853;
    wire N__1848;
    wire N__1845;
    wire N__1842;
    wire N__1835;
    wire N__1832;
    wire N__1829;
    wire N__1826;
    wire N__1823;
    wire N__1820;
    wire N__1817;
    wire N__1814;
    wire N__1811;
    wire N__1808;
    wire N__1805;
    wire N__1802;
    wire N__1801;
    wire N__1800;
    wire N__1799;
    wire N__1790;
    wire N__1787;
    wire N__1784;
    wire N__1781;
    wire N__1780;
    wire N__1777;
    wire N__1774;
    wire N__1769;
    wire N__1768;
    wire N__1765;
    wire N__1762;
    wire N__1757;
    wire N__1754;
    wire N__1753;
    wire N__1750;
    wire N__1747;
    wire N__1742;
    wire N__1741;
    wire N__1738;
    wire N__1735;
    wire N__1730;
    wire N__1727;
    wire N__1724;
    wire N__1723;
    wire N__1720;
    wire N__1717;
    wire N__1714;
    wire N__1709;
    wire N__1708;
    wire N__1705;
    wire N__1702;
    wire N__1697;
    wire N__1696;
    wire N__1693;
    wire N__1690;
    wire N__1685;
    wire N__1684;
    wire N__1681;
    wire N__1678;
    wire N__1673;
    wire N__1670;
    wire N__1667;
    wire N__1664;
    wire N__1661;
    wire N__1658;
    wire N__1655;
    wire N__1652;
    wire N__1649;
    wire N__1646;
    wire N__1643;
    wire N__1640;
    wire N__1637;
    wire N__1634;
    wire N__1633;
    wire N__1628;
    wire N__1625;
    wire N__1624;
    wire N__1619;
    wire N__1616;
    wire N__1613;
    wire N__1612;
    wire N__1607;
    wire N__1604;
    wire N__1603;
    wire N__1598;
    wire N__1595;
    wire N__1594;
    wire N__1593;
    wire N__1592;
    wire N__1589;
    wire N__1582;
    wire N__1577;
    wire N__1576;
    wire N__1573;
    wire N__1570;
    wire N__1569;
    wire N__1566;
    wire N__1561;
    wire N__1556;
    wire N__1555;
    wire N__1552;
    wire N__1549;
    wire N__1544;
    wire N__1541;
    wire N__1540;
    wire N__1537;
    wire N__1534;
    wire N__1531;
    wire N__1526;
    wire N__1523;
    wire N__1522;
    wire N__1519;
    wire N__1516;
    wire N__1511;
    wire N__1508;
    wire N__1505;
    wire N__1502;
    wire N__1499;
    wire N__1496;
    wire N__1493;
    wire N__1490;
    wire N__1487;
    wire N__1484;
    wire N__1481;
    wire N__1478;
    wire N__1475;
    wire N__1472;
    wire N__1469;
    wire N__1466;
    wire N__1463;
    wire N__1460;
    wire N__1457;
    wire N__1454;
    wire N__1451;
    wire N__1448;
    wire N__1445;
    wire N__1442;
    wire N__1439;
    wire N__1436;
    wire N__1433;
    wire N__1430;
    wire N__1427;
    wire N__1424;
    wire VCCG0;
    wire GNDG0;
    wire \Debounce_Sw1.un9_r_count_10_cascade_ ;
    wire \Debounce_Sw1.un1_r_Count_1lt11_0_cascade_ ;
    wire \Debounce_Sw1.un1_r_Count_1lto11_1 ;
    wire \Debounce_Sw1.un1_r_Count_1lt17_cascade_ ;
    wire \Debounce_Sw1.un1_r_Count_1lto17_2 ;
    wire \Debounce_Sw1.r_count15_i ;
    wire bfn_4_7_0_;
    wire \Count_And_Toggle.un2_r_counter_cry_1 ;
    wire \Count_And_Toggle.un2_r_counter_cry_2 ;
    wire \Count_And_Toggle.un2_r_counter_cry_3 ;
    wire \Count_And_Toggle.un2_r_counter_cry_4 ;
    wire \Count_And_Toggle.un2_r_counter_cry_5 ;
    wire \Count_And_Toggle.un2_r_counter_cry_6 ;
    wire \Count_And_Toggle.un2_r_counter_cry_7 ;
    wire \Count_And_Toggle.un2_r_counter_cry_8 ;
    wire bfn_4_8_0_;
    wire \Count_And_Toggle.un2_r_counter_cry_9 ;
    wire \Count_And_Toggle.un2_r_counter_cry_10 ;
    wire \Count_And_Toggle.un2_r_counter_cry_11 ;
    wire \Count_And_Toggle.un2_r_counter_cry_12 ;
    wire \Count_And_Toggle.un2_r_counter_cry_13 ;
    wire \Count_And_Toggle.un2_r_counter_cry_14 ;
    wire \Count_And_Toggle.un2_r_counter_cry_15 ;
    wire \Count_And_Toggle.un2_r_counter_cry_16 ;
    wire bfn_4_9_0_;
    wire \Count_And_Toggle.un2_r_counter_cry_17 ;
    wire \Count_And_Toggle.un2_r_counter_cry_18 ;
    wire \Count_And_Toggle.un2_r_counter_cry_19 ;
    wire \Count_And_Toggle.un2_r_counter_cry_20 ;
    wire \Count_And_Toggle.un2_r_counter_cry_21 ;
    wire \Count_And_Toggle.r_Counter_RNO_0Z0Z_22_cascade_ ;
    wire \Count_And_Toggle.r_CounterZ0Z_17 ;
    wire \Count_And_Toggle.r_CounterZ0Z_22 ;
    wire \Count_And_Toggle.r_CounterZ0Z_21 ;
    wire \Count_And_Toggle.r_CounterZ0Z_20 ;
    wire \Debounce_Sw1.r_CountZ0Z_0 ;
    wire \Debounce_Sw1.r_CountZ0Z_1 ;
    wire bfn_5_5_0_;
    wire \Debounce_Sw1.r_CountZ0Z_2 ;
    wire \Debounce_Sw1.un2_r_count_cry_1 ;
    wire \Debounce_Sw1.r_CountZ0Z_3 ;
    wire \Debounce_Sw1.un2_r_count_cry_2 ;
    wire \Debounce_Sw1.r_CountZ0Z_4 ;
    wire \Debounce_Sw1.un2_r_count_cry_3 ;
    wire \Debounce_Sw1.r_CountZ0Z_5 ;
    wire \Debounce_Sw1.un2_r_count_cry_4 ;
    wire \Debounce_Sw1.un2_r_count_cry_5 ;
    wire \Debounce_Sw1.un2_r_count_cry_6 ;
    wire \Debounce_Sw1.un2_r_count_cry_7 ;
    wire \Debounce_Sw1.un2_r_count_cry_8 ;
    wire bfn_5_6_0_;
    wire \Debounce_Sw1.un2_r_count_cry_9 ;
    wire \Debounce_Sw1.un2_r_count_cry_10 ;
    wire \Debounce_Sw1.un2_r_count_cry_11 ;
    wire \Debounce_Sw1.un2_r_count_cry_12 ;
    wire \Debounce_Sw1.un2_r_count_cry_13 ;
    wire \Debounce_Sw1.un2_r_count_cry_14 ;
    wire \Debounce_Sw1.un2_r_count_cry_15 ;
    wire \Debounce_Sw1.un2_r_count_cry_16 ;
    wire bfn_5_7_0_;
    wire \Debounce_Sw1.r_count15_i_g ;
    wire \Count_And_Toggle.r_CounterZ0Z_12 ;
    wire \Count_And_Toggle.r_CounterZ0Z_10 ;
    wire \Count_And_Toggle.r_CounterZ0Z_13 ;
    wire \Count_And_Toggle.r_CounterZ0Z_7 ;
    wire \Count_And_Toggle.r_Counter_RNO_0Z0Z_8 ;
    wire \Count_And_Toggle.r_CounterZ0Z_8 ;
    wire \Count_And_Toggle.r_CounterZ0Z_5 ;
    wire \Count_And_Toggle.r_CounterZ0Z_4 ;
    wire \Count_And_Toggle.r_Counter_RNO_0Z0Z_11 ;
    wire \Count_And_Toggle.r_CounterZ0Z_3 ;
    wire \Count_And_Toggle.r_CounterZ0Z_2 ;
    wire \Count_And_Toggle.r_CounterZ0Z_1 ;
    wire \Count_And_Toggle.r_Counter_RNO_0Z0Z_6 ;
    wire \Count_And_Toggle.r_CounterZ0Z_6 ;
    wire \Count_And_Toggle.r_Counter_RNO_0Z0Z_19 ;
    wire \Count_And_Toggle.r_CounterZ0Z_19 ;
    wire \Count_And_Toggle.r_CounterZ0Z_11 ;
    wire \Count_And_Toggle.un4_i_enable_15_cascade_ ;
    wire \Count_And_Toggle.r_Counter_RNO_0Z0Z_18 ;
    wire \Count_And_Toggle.r_CounterZ0Z_18 ;
    wire \Count_And_Toggle.r_CounterZ0Z_15 ;
    wire \Count_And_Toggle.r_CounterZ0Z_16 ;
    wire \Count_And_Toggle.r_CounterZ0Z_0 ;
    wire \Count_And_Toggle.un4_i_enable_14 ;
    wire \Count_And_Toggle.un4_i_enable_12 ;
    wire \Count_And_Toggle.un4_i_enable_11_cascade_ ;
    wire \Count_And_Toggle.un4_i_enable_13 ;
    wire \Count_And_Toggle.un4_i_enable_20_cascade_ ;
    wire \Count_And_Toggle.r_Counter_RNO_0Z0Z_14 ;
    wire \Count_And_Toggle.r_CounterZ0Z_14 ;
    wire \Debounce_Sw1.r_CountZ0Z_8 ;
    wire \Debounce_Sw1.r_CountZ0Z_6 ;
    wire \Debounce_Sw1.un9_r_count_9 ;
    wire \Debounce_Sw1.r_CountZ0Z_12 ;
    wire \Debounce_Sw1.r_CountZ0Z_14 ;
    wire \Debounce_Sw1.r_CountZ0Z_15 ;
    wire \Debounce_Sw1.r_CountZ0Z_7 ;
    wire \Debounce_Sw1.un9_r_count_10 ;
    wire \Debounce_Sw1.r_CountZ0Z_9 ;
    wire \Debounce_Sw1.un9_r_count_5_cascade_ ;
    wire \Debounce_Sw1.r_CountZ0Z_10 ;
    wire \Debounce_Sw1.un9_r_count_9_0 ;
    wire i_Switch_1_c;
    wire \Debounce_Sw1.un9_r_count_10_0_cascade_ ;
    wire \Debounce_Sw1.r_CountZ0Z_16 ;
    wire \Debounce_Sw1.r_CountZ0Z_13 ;
    wire \Debounce_Sw1.r_CountZ0Z_17 ;
    wire \Debounce_Sw1.r_CountZ0Z_11 ;
    wire \Debounce_Sw1.un9_r_count_6 ;
    wire \Count_And_Toggle.r_Counter_RNO_0Z0Z_9 ;
    wire \Count_And_Toggle.r_CounterZ0Z_9 ;
    wire \Count_And_Toggle.un4_i_enable_16 ;
    wire \Count_And_Toggle.un4_i_enable_15 ;
    wire \Count_And_Toggle.un4_i_enable_20 ;
    wire \Debounce_Sw2.un9_r_count_10_cascade_ ;
    wire \Debounce_Sw2.N_23_cascade_ ;
    wire i_Switch_2_c;
    wire \Debounce_Sw2.N_16_cascade_ ;
    wire \Debounce_Sw2.N_9 ;
    wire \Debounce_Sw2.un9_r_count_10 ;
    wire \Debounce_Sw2.r_State_e_0_RNOZ0 ;
    wire \Debounce_Sw2.N_10 ;
    wire \Debounce_Sw2.un9_r_count_0_a3_2 ;
    wire \Debounce_Sw2.N_22_3 ;
    wire \Debounce_Sw2.N_13 ;
    wire \Debounce_Sw2.r_CountZ0Z_0 ;
    wire \Debounce_Sw2.r_CountZ0Z_1 ;
    wire bfn_8_9_0_;
    wire \Debounce_Sw2.r_CountZ0Z_2 ;
    wire \Debounce_Sw2.un2_r_count_cry_1 ;
    wire \Debounce_Sw2.r_CountZ0Z_3 ;
    wire \Debounce_Sw2.un2_r_count_cry_2 ;
    wire \Debounce_Sw2.r_CountZ0Z_4 ;
    wire \Debounce_Sw2.un2_r_count_cry_3 ;
    wire \Debounce_Sw2.r_CountZ0Z_5 ;
    wire \Debounce_Sw2.un2_r_count_cry_4 ;
    wire \Debounce_Sw2.r_CountZ0Z_6 ;
    wire \Debounce_Sw2.un2_r_count_cry_5 ;
    wire \Debounce_Sw2.r_CountZ0Z_7 ;
    wire \Debounce_Sw2.un2_r_count_cry_6 ;
    wire \Debounce_Sw2.r_CountZ0Z_8 ;
    wire \Debounce_Sw2.un2_r_count_cry_7 ;
    wire \Debounce_Sw2.un2_r_count_cry_8 ;
    wire \Debounce_Sw2.r_CountZ0Z_9 ;
    wire bfn_8_10_0_;
    wire \Debounce_Sw2.r_CountZ0Z_10 ;
    wire \Debounce_Sw2.un2_r_count_cry_9 ;
    wire \Debounce_Sw2.r_CountZ0Z_11 ;
    wire \Debounce_Sw2.un2_r_count_cry_10 ;
    wire \Debounce_Sw2.r_CountZ0Z_12 ;
    wire \Debounce_Sw2.un2_r_count_cry_11 ;
    wire \Debounce_Sw2.r_CountZ0Z_13 ;
    wire \Debounce_Sw2.un2_r_count_cry_12 ;
    wire \Debounce_Sw2.r_CountZ0Z_14 ;
    wire \Debounce_Sw2.un2_r_count_cry_13 ;
    wire \Debounce_Sw2.r_CountZ0Z_15 ;
    wire \Debounce_Sw2.un2_r_count_cry_14 ;
    wire \Debounce_Sw2.r_CountZ0Z_16 ;
    wire \Debounce_Sw2.un2_r_count_cry_15 ;
    wire \Debounce_Sw2.un2_r_count_cry_16 ;
    wire bfn_8_11_0_;
    wire \Debounce_Sw2.r_CountZ0Z_17 ;
    wire i_Clk_c_g;
    wire \Debounce_Sw2.N_9_g ;
    wire o_LED_2_c;
    wire o_LED_3_c;
    wire o_LED_1_c;
    wire w_Switch_1;
    wire w_Toggle;
    wire w_Switch_2;
    wire o_LED_4_c;
    wire _gnd_net_;

    PRE_IO_GBUF i_Clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__3210),
            .GLOBALBUFFEROUTPUT(i_Clk_c_g));
    IO_PAD i_Clk_ibuf_gb_io_iopad (
            .OE(N__3212),
            .DIN(N__3211),
            .DOUT(N__3210),
            .PACKAGEPIN(i_Clk));
    defparam i_Clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam i_Clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Clk_ibuf_gb_io_preio (
            .PADOEN(N__3212),
            .PADOUT(N__3211),
            .PADIN(N__3210),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_1_obuf_iopad (
            .OE(N__3201),
            .DIN(N__3200),
            .DOUT(N__3199),
            .PACKAGEPIN(o_LED_1));
    defparam o_LED_1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_1_obuf_preio (
            .PADOEN(N__3201),
            .PADOUT(N__3200),
            .PADIN(N__3199),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2999),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_1_ibuf_iopad (
            .OE(N__3192),
            .DIN(N__3191),
            .DOUT(N__3190),
            .PACKAGEPIN(i_Switch_1));
    defparam i_Switch_1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_1_ibuf_preio (
            .PADOEN(N__3192),
            .PADOUT(N__3191),
            .PADIN(N__3190),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_2_obuf_iopad (
            .OE(N__3183),
            .DIN(N__3182),
            .DOUT(N__3181),
            .PACKAGEPIN(o_LED_2));
    defparam o_LED_2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_2_obuf_preio (
            .PADOEN(N__3183),
            .PADOUT(N__3182),
            .PADIN(N__3181),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3011),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_2_ibuf_iopad (
            .OE(N__3174),
            .DIN(N__3173),
            .DOUT(N__3172),
            .PACKAGEPIN(i_Switch_2));
    defparam i_Switch_2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_2_ibuf_preio (
            .PADOEN(N__3174),
            .PADOUT(N__3173),
            .PADIN(N__3172),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_3_obuf_iopad (
            .OE(N__3165),
            .DIN(N__3164),
            .DOUT(N__3163),
            .PACKAGEPIN(o_LED_3));
    defparam o_LED_3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_3_obuf_preio (
            .PADOEN(N__3165),
            .PADOUT(N__3164),
            .PADIN(N__3163),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3005),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_4_obuf_iopad (
            .OE(N__3156),
            .DIN(N__3155),
            .DOUT(N__3154),
            .PACKAGEPIN(o_LED_4));
    defparam o_LED_4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_4_obuf_preio (
            .PADOEN(N__3156),
            .PADOUT(N__3155),
            .PADIN(N__3154),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2882),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__696 (
            .O(N__3137),
            .I(N__3133));
    InMux I__695 (
            .O(N__3136),
            .I(N__3130));
    LocalMux I__694 (
            .O(N__3133),
            .I(\Debounce_Sw2.r_CountZ0Z_15 ));
    LocalMux I__693 (
            .O(N__3130),
            .I(\Debounce_Sw2.r_CountZ0Z_15 ));
    InMux I__692 (
            .O(N__3125),
            .I(\Debounce_Sw2.un2_r_count_cry_14 ));
    InMux I__691 (
            .O(N__3122),
            .I(N__3118));
    InMux I__690 (
            .O(N__3121),
            .I(N__3115));
    LocalMux I__689 (
            .O(N__3118),
            .I(\Debounce_Sw2.r_CountZ0Z_16 ));
    LocalMux I__688 (
            .O(N__3115),
            .I(\Debounce_Sw2.r_CountZ0Z_16 ));
    InMux I__687 (
            .O(N__3110),
            .I(\Debounce_Sw2.un2_r_count_cry_15 ));
    InMux I__686 (
            .O(N__3107),
            .I(bfn_8_11_0_));
    CascadeMux I__685 (
            .O(N__3104),
            .I(N__3101));
    InMux I__684 (
            .O(N__3101),
            .I(N__3097));
    InMux I__683 (
            .O(N__3100),
            .I(N__3094));
    LocalMux I__682 (
            .O(N__3097),
            .I(N__3091));
    LocalMux I__681 (
            .O(N__3094),
            .I(\Debounce_Sw2.r_CountZ0Z_17 ));
    Odrv4 I__680 (
            .O(N__3091),
            .I(\Debounce_Sw2.r_CountZ0Z_17 ));
    ClkMux I__679 (
            .O(N__3086),
            .I(N__3035));
    ClkMux I__678 (
            .O(N__3085),
            .I(N__3035));
    ClkMux I__677 (
            .O(N__3084),
            .I(N__3035));
    ClkMux I__676 (
            .O(N__3083),
            .I(N__3035));
    ClkMux I__675 (
            .O(N__3082),
            .I(N__3035));
    ClkMux I__674 (
            .O(N__3081),
            .I(N__3035));
    ClkMux I__673 (
            .O(N__3080),
            .I(N__3035));
    ClkMux I__672 (
            .O(N__3079),
            .I(N__3035));
    ClkMux I__671 (
            .O(N__3078),
            .I(N__3035));
    ClkMux I__670 (
            .O(N__3077),
            .I(N__3035));
    ClkMux I__669 (
            .O(N__3076),
            .I(N__3035));
    ClkMux I__668 (
            .O(N__3075),
            .I(N__3035));
    ClkMux I__667 (
            .O(N__3074),
            .I(N__3035));
    ClkMux I__666 (
            .O(N__3073),
            .I(N__3035));
    ClkMux I__665 (
            .O(N__3072),
            .I(N__3035));
    ClkMux I__664 (
            .O(N__3071),
            .I(N__3035));
    ClkMux I__663 (
            .O(N__3070),
            .I(N__3035));
    GlobalMux I__662 (
            .O(N__3035),
            .I(N__3032));
    gio2CtrlBuf I__661 (
            .O(N__3032),
            .I(i_Clk_c_g));
    SRMux I__660 (
            .O(N__3029),
            .I(N__3017));
    SRMux I__659 (
            .O(N__3028),
            .I(N__3017));
    SRMux I__658 (
            .O(N__3027),
            .I(N__3017));
    SRMux I__657 (
            .O(N__3026),
            .I(N__3017));
    GlobalMux I__656 (
            .O(N__3017),
            .I(N__3014));
    gio2CtrlBuf I__655 (
            .O(N__3014),
            .I(\Debounce_Sw2.N_9_g ));
    IoInMux I__654 (
            .O(N__3011),
            .I(N__3008));
    LocalMux I__653 (
            .O(N__3008),
            .I(o_LED_2_c));
    IoInMux I__652 (
            .O(N__3005),
            .I(N__3002));
    LocalMux I__651 (
            .O(N__3002),
            .I(o_LED_3_c));
    IoInMux I__650 (
            .O(N__2999),
            .I(N__2996));
    LocalMux I__649 (
            .O(N__2996),
            .I(o_LED_1_c));
    InMux I__648 (
            .O(N__2993),
            .I(N__2987));
    InMux I__647 (
            .O(N__2992),
            .I(N__2980));
    InMux I__646 (
            .O(N__2991),
            .I(N__2980));
    InMux I__645 (
            .O(N__2990),
            .I(N__2980));
    LocalMux I__644 (
            .O(N__2987),
            .I(N__2975));
    LocalMux I__643 (
            .O(N__2980),
            .I(N__2975));
    Span4Mux_v I__642 (
            .O(N__2975),
            .I(N__2970));
    InMux I__641 (
            .O(N__2974),
            .I(N__2967));
    InMux I__640 (
            .O(N__2973),
            .I(N__2964));
    Span4Mux_h I__639 (
            .O(N__2970),
            .I(N__2959));
    LocalMux I__638 (
            .O(N__2967),
            .I(N__2959));
    LocalMux I__637 (
            .O(N__2964),
            .I(w_Switch_1));
    Odrv4 I__636 (
            .O(N__2959),
            .I(w_Switch_1));
    InMux I__635 (
            .O(N__2954),
            .I(N__2944));
    InMux I__634 (
            .O(N__2953),
            .I(N__2944));
    InMux I__633 (
            .O(N__2952),
            .I(N__2944));
    InMux I__632 (
            .O(N__2951),
            .I(N__2941));
    LocalMux I__631 (
            .O(N__2944),
            .I(N__2936));
    LocalMux I__630 (
            .O(N__2941),
            .I(N__2936));
    Span4Mux_v I__629 (
            .O(N__2936),
            .I(N__2932));
    CascadeMux I__628 (
            .O(N__2935),
            .I(N__2929));
    Span4Mux_h I__627 (
            .O(N__2932),
            .I(N__2926));
    InMux I__626 (
            .O(N__2929),
            .I(N__2923));
    Odrv4 I__625 (
            .O(N__2926),
            .I(w_Toggle));
    LocalMux I__624 (
            .O(N__2923),
            .I(w_Toggle));
    CascadeMux I__623 (
            .O(N__2918),
            .I(N__2914));
    InMux I__622 (
            .O(N__2917),
            .I(N__2905));
    InMux I__621 (
            .O(N__2914),
            .I(N__2905));
    InMux I__620 (
            .O(N__2913),
            .I(N__2905));
    InMux I__619 (
            .O(N__2912),
            .I(N__2902));
    LocalMux I__618 (
            .O(N__2905),
            .I(N__2897));
    LocalMux I__617 (
            .O(N__2902),
            .I(N__2897));
    Span4Mux_v I__616 (
            .O(N__2897),
            .I(N__2894));
    Span4Mux_h I__615 (
            .O(N__2894),
            .I(N__2890));
    InMux I__614 (
            .O(N__2893),
            .I(N__2887));
    Odrv4 I__613 (
            .O(N__2890),
            .I(w_Switch_2));
    LocalMux I__612 (
            .O(N__2887),
            .I(w_Switch_2));
    IoInMux I__611 (
            .O(N__2882),
            .I(N__2879));
    LocalMux I__610 (
            .O(N__2879),
            .I(o_LED_4_c));
    InMux I__609 (
            .O(N__2876),
            .I(N__2872));
    InMux I__608 (
            .O(N__2875),
            .I(N__2869));
    LocalMux I__607 (
            .O(N__2872),
            .I(\Debounce_Sw2.r_CountZ0Z_6 ));
    LocalMux I__606 (
            .O(N__2869),
            .I(\Debounce_Sw2.r_CountZ0Z_6 ));
    InMux I__605 (
            .O(N__2864),
            .I(\Debounce_Sw2.un2_r_count_cry_5 ));
    CascadeMux I__604 (
            .O(N__2861),
            .I(N__2857));
    InMux I__603 (
            .O(N__2860),
            .I(N__2853));
    InMux I__602 (
            .O(N__2857),
            .I(N__2850));
    InMux I__601 (
            .O(N__2856),
            .I(N__2847));
    LocalMux I__600 (
            .O(N__2853),
            .I(\Debounce_Sw2.r_CountZ0Z_7 ));
    LocalMux I__599 (
            .O(N__2850),
            .I(\Debounce_Sw2.r_CountZ0Z_7 ));
    LocalMux I__598 (
            .O(N__2847),
            .I(\Debounce_Sw2.r_CountZ0Z_7 ));
    InMux I__597 (
            .O(N__2840),
            .I(\Debounce_Sw2.un2_r_count_cry_6 ));
    InMux I__596 (
            .O(N__2837),
            .I(N__2833));
    InMux I__595 (
            .O(N__2836),
            .I(N__2830));
    LocalMux I__594 (
            .O(N__2833),
            .I(\Debounce_Sw2.r_CountZ0Z_8 ));
    LocalMux I__593 (
            .O(N__2830),
            .I(\Debounce_Sw2.r_CountZ0Z_8 ));
    InMux I__592 (
            .O(N__2825),
            .I(\Debounce_Sw2.un2_r_count_cry_7 ));
    InMux I__591 (
            .O(N__2822),
            .I(N__2818));
    InMux I__590 (
            .O(N__2821),
            .I(N__2815));
    LocalMux I__589 (
            .O(N__2818),
            .I(\Debounce_Sw2.r_CountZ0Z_9 ));
    LocalMux I__588 (
            .O(N__2815),
            .I(\Debounce_Sw2.r_CountZ0Z_9 ));
    InMux I__587 (
            .O(N__2810),
            .I(bfn_8_10_0_));
    InMux I__586 (
            .O(N__2807),
            .I(N__2803));
    InMux I__585 (
            .O(N__2806),
            .I(N__2800));
    LocalMux I__584 (
            .O(N__2803),
            .I(\Debounce_Sw2.r_CountZ0Z_10 ));
    LocalMux I__583 (
            .O(N__2800),
            .I(\Debounce_Sw2.r_CountZ0Z_10 ));
    InMux I__582 (
            .O(N__2795),
            .I(\Debounce_Sw2.un2_r_count_cry_9 ));
    CascadeMux I__581 (
            .O(N__2792),
            .I(N__2788));
    InMux I__580 (
            .O(N__2791),
            .I(N__2785));
    InMux I__579 (
            .O(N__2788),
            .I(N__2782));
    LocalMux I__578 (
            .O(N__2785),
            .I(\Debounce_Sw2.r_CountZ0Z_11 ));
    LocalMux I__577 (
            .O(N__2782),
            .I(\Debounce_Sw2.r_CountZ0Z_11 ));
    InMux I__576 (
            .O(N__2777),
            .I(\Debounce_Sw2.un2_r_count_cry_10 ));
    InMux I__575 (
            .O(N__2774),
            .I(N__2769));
    InMux I__574 (
            .O(N__2773),
            .I(N__2764));
    InMux I__573 (
            .O(N__2772),
            .I(N__2764));
    LocalMux I__572 (
            .O(N__2769),
            .I(\Debounce_Sw2.r_CountZ0Z_12 ));
    LocalMux I__571 (
            .O(N__2764),
            .I(\Debounce_Sw2.r_CountZ0Z_12 ));
    InMux I__570 (
            .O(N__2759),
            .I(\Debounce_Sw2.un2_r_count_cry_11 ));
    InMux I__569 (
            .O(N__2756),
            .I(N__2751));
    InMux I__568 (
            .O(N__2755),
            .I(N__2748));
    InMux I__567 (
            .O(N__2754),
            .I(N__2745));
    LocalMux I__566 (
            .O(N__2751),
            .I(\Debounce_Sw2.r_CountZ0Z_13 ));
    LocalMux I__565 (
            .O(N__2748),
            .I(\Debounce_Sw2.r_CountZ0Z_13 ));
    LocalMux I__564 (
            .O(N__2745),
            .I(\Debounce_Sw2.r_CountZ0Z_13 ));
    InMux I__563 (
            .O(N__2738),
            .I(\Debounce_Sw2.un2_r_count_cry_12 ));
    InMux I__562 (
            .O(N__2735),
            .I(N__2731));
    InMux I__561 (
            .O(N__2734),
            .I(N__2728));
    LocalMux I__560 (
            .O(N__2731),
            .I(\Debounce_Sw2.r_CountZ0Z_14 ));
    LocalMux I__559 (
            .O(N__2728),
            .I(\Debounce_Sw2.r_CountZ0Z_14 ));
    InMux I__558 (
            .O(N__2723),
            .I(\Debounce_Sw2.un2_r_count_cry_13 ));
    InMux I__557 (
            .O(N__2720),
            .I(N__2716));
    InMux I__556 (
            .O(N__2719),
            .I(N__2713));
    LocalMux I__555 (
            .O(N__2716),
            .I(\Debounce_Sw2.N_10 ));
    LocalMux I__554 (
            .O(N__2713),
            .I(\Debounce_Sw2.N_10 ));
    InMux I__553 (
            .O(N__2708),
            .I(N__2705));
    LocalMux I__552 (
            .O(N__2705),
            .I(\Debounce_Sw2.un9_r_count_0_a3_2 ));
    InMux I__551 (
            .O(N__2702),
            .I(N__2696));
    InMux I__550 (
            .O(N__2701),
            .I(N__2696));
    LocalMux I__549 (
            .O(N__2696),
            .I(\Debounce_Sw2.N_22_3 ));
    InMux I__548 (
            .O(N__2693),
            .I(N__2687));
    InMux I__547 (
            .O(N__2692),
            .I(N__2687));
    LocalMux I__546 (
            .O(N__2687),
            .I(\Debounce_Sw2.N_13 ));
    InMux I__545 (
            .O(N__2684),
            .I(N__2676));
    InMux I__544 (
            .O(N__2683),
            .I(N__2676));
    InMux I__543 (
            .O(N__2682),
            .I(N__2673));
    InMux I__542 (
            .O(N__2681),
            .I(N__2670));
    LocalMux I__541 (
            .O(N__2676),
            .I(\Debounce_Sw2.r_CountZ0Z_0 ));
    LocalMux I__540 (
            .O(N__2673),
            .I(\Debounce_Sw2.r_CountZ0Z_0 ));
    LocalMux I__539 (
            .O(N__2670),
            .I(\Debounce_Sw2.r_CountZ0Z_0 ));
    CascadeMux I__538 (
            .O(N__2663),
            .I(N__2659));
    InMux I__537 (
            .O(N__2662),
            .I(N__2655));
    InMux I__536 (
            .O(N__2659),
            .I(N__2652));
    InMux I__535 (
            .O(N__2658),
            .I(N__2649));
    LocalMux I__534 (
            .O(N__2655),
            .I(\Debounce_Sw2.r_CountZ0Z_1 ));
    LocalMux I__533 (
            .O(N__2652),
            .I(\Debounce_Sw2.r_CountZ0Z_1 ));
    LocalMux I__532 (
            .O(N__2649),
            .I(\Debounce_Sw2.r_CountZ0Z_1 ));
    CascadeMux I__531 (
            .O(N__2642),
            .I(N__2639));
    InMux I__530 (
            .O(N__2639),
            .I(N__2635));
    InMux I__529 (
            .O(N__2638),
            .I(N__2632));
    LocalMux I__528 (
            .O(N__2635),
            .I(N__2629));
    LocalMux I__527 (
            .O(N__2632),
            .I(\Debounce_Sw2.r_CountZ0Z_2 ));
    Odrv4 I__526 (
            .O(N__2629),
            .I(\Debounce_Sw2.r_CountZ0Z_2 ));
    InMux I__525 (
            .O(N__2624),
            .I(\Debounce_Sw2.un2_r_count_cry_1 ));
    InMux I__524 (
            .O(N__2621),
            .I(N__2617));
    InMux I__523 (
            .O(N__2620),
            .I(N__2614));
    LocalMux I__522 (
            .O(N__2617),
            .I(\Debounce_Sw2.r_CountZ0Z_3 ));
    LocalMux I__521 (
            .O(N__2614),
            .I(\Debounce_Sw2.r_CountZ0Z_3 ));
    InMux I__520 (
            .O(N__2609),
            .I(\Debounce_Sw2.un2_r_count_cry_2 ));
    InMux I__519 (
            .O(N__2606),
            .I(N__2602));
    InMux I__518 (
            .O(N__2605),
            .I(N__2599));
    LocalMux I__517 (
            .O(N__2602),
            .I(\Debounce_Sw2.r_CountZ0Z_4 ));
    LocalMux I__516 (
            .O(N__2599),
            .I(\Debounce_Sw2.r_CountZ0Z_4 ));
    InMux I__515 (
            .O(N__2594),
            .I(\Debounce_Sw2.un2_r_count_cry_3 ));
    InMux I__514 (
            .O(N__2591),
            .I(N__2587));
    InMux I__513 (
            .O(N__2590),
            .I(N__2584));
    LocalMux I__512 (
            .O(N__2587),
            .I(N__2581));
    LocalMux I__511 (
            .O(N__2584),
            .I(\Debounce_Sw2.r_CountZ0Z_5 ));
    Odrv4 I__510 (
            .O(N__2581),
            .I(\Debounce_Sw2.r_CountZ0Z_5 ));
    InMux I__509 (
            .O(N__2576),
            .I(\Debounce_Sw2.un2_r_count_cry_4 ));
    InMux I__508 (
            .O(N__2573),
            .I(N__2563));
    InMux I__507 (
            .O(N__2572),
            .I(N__2560));
    InMux I__506 (
            .O(N__2571),
            .I(N__2553));
    InMux I__505 (
            .O(N__2570),
            .I(N__2553));
    InMux I__504 (
            .O(N__2569),
            .I(N__2553));
    InMux I__503 (
            .O(N__2568),
            .I(N__2550));
    InMux I__502 (
            .O(N__2567),
            .I(N__2545));
    InMux I__501 (
            .O(N__2566),
            .I(N__2545));
    LocalMux I__500 (
            .O(N__2563),
            .I(\Count_And_Toggle.un4_i_enable_20 ));
    LocalMux I__499 (
            .O(N__2560),
            .I(\Count_And_Toggle.un4_i_enable_20 ));
    LocalMux I__498 (
            .O(N__2553),
            .I(\Count_And_Toggle.un4_i_enable_20 ));
    LocalMux I__497 (
            .O(N__2550),
            .I(\Count_And_Toggle.un4_i_enable_20 ));
    LocalMux I__496 (
            .O(N__2545),
            .I(\Count_And_Toggle.un4_i_enable_20 ));
    CascadeMux I__495 (
            .O(N__2534),
            .I(\Debounce_Sw2.un9_r_count_10_cascade_ ));
    CascadeMux I__494 (
            .O(N__2531),
            .I(\Debounce_Sw2.N_23_cascade_ ));
    InMux I__493 (
            .O(N__2528),
            .I(N__2525));
    LocalMux I__492 (
            .O(N__2525),
            .I(N__2521));
    InMux I__491 (
            .O(N__2524),
            .I(N__2518));
    Span4Mux_v I__490 (
            .O(N__2521),
            .I(N__2515));
    LocalMux I__489 (
            .O(N__2518),
            .I(N__2512));
    Span4Mux_h I__488 (
            .O(N__2515),
            .I(N__2509));
    Span12Mux_v I__487 (
            .O(N__2512),
            .I(N__2506));
    Span4Mux_v I__486 (
            .O(N__2509),
            .I(N__2503));
    Odrv12 I__485 (
            .O(N__2506),
            .I(i_Switch_2_c));
    Odrv4 I__484 (
            .O(N__2503),
            .I(i_Switch_2_c));
    CascadeMux I__483 (
            .O(N__2498),
            .I(\Debounce_Sw2.N_16_cascade_ ));
    IoInMux I__482 (
            .O(N__2495),
            .I(N__2492));
    LocalMux I__481 (
            .O(N__2492),
            .I(N__2489));
    Span12Mux_s7_v I__480 (
            .O(N__2489),
            .I(N__2486));
    Odrv12 I__479 (
            .O(N__2486),
            .I(\Debounce_Sw2.N_9 ));
    CascadeMux I__478 (
            .O(N__2483),
            .I(N__2480));
    InMux I__477 (
            .O(N__2480),
            .I(N__2477));
    LocalMux I__476 (
            .O(N__2477),
            .I(\Debounce_Sw2.un9_r_count_10 ));
    CEMux I__475 (
            .O(N__2474),
            .I(N__2471));
    LocalMux I__474 (
            .O(N__2471),
            .I(N__2468));
    Odrv4 I__473 (
            .O(N__2468),
            .I(\Debounce_Sw2.r_State_e_0_RNOZ0 ));
    CascadeMux I__472 (
            .O(N__2465),
            .I(\Count_And_Toggle.un4_i_enable_20_cascade_ ));
    InMux I__471 (
            .O(N__2462),
            .I(N__2459));
    LocalMux I__470 (
            .O(N__2459),
            .I(\Count_And_Toggle.r_Counter_RNO_0Z0Z_14 ));
    InMux I__469 (
            .O(N__2456),
            .I(N__2452));
    InMux I__468 (
            .O(N__2455),
            .I(N__2449));
    LocalMux I__467 (
            .O(N__2452),
            .I(\Count_And_Toggle.r_CounterZ0Z_14 ));
    LocalMux I__466 (
            .O(N__2449),
            .I(\Count_And_Toggle.r_CounterZ0Z_14 ));
    InMux I__465 (
            .O(N__2444),
            .I(N__2439));
    InMux I__464 (
            .O(N__2443),
            .I(N__2436));
    InMux I__463 (
            .O(N__2442),
            .I(N__2433));
    LocalMux I__462 (
            .O(N__2439),
            .I(\Debounce_Sw1.r_CountZ0Z_8 ));
    LocalMux I__461 (
            .O(N__2436),
            .I(\Debounce_Sw1.r_CountZ0Z_8 ));
    LocalMux I__460 (
            .O(N__2433),
            .I(\Debounce_Sw1.r_CountZ0Z_8 ));
    CascadeMux I__459 (
            .O(N__2426),
            .I(N__2423));
    InMux I__458 (
            .O(N__2423),
            .I(N__2418));
    InMux I__457 (
            .O(N__2422),
            .I(N__2415));
    InMux I__456 (
            .O(N__2421),
            .I(N__2412));
    LocalMux I__455 (
            .O(N__2418),
            .I(\Debounce_Sw1.r_CountZ0Z_6 ));
    LocalMux I__454 (
            .O(N__2415),
            .I(\Debounce_Sw1.r_CountZ0Z_6 ));
    LocalMux I__453 (
            .O(N__2412),
            .I(\Debounce_Sw1.r_CountZ0Z_6 ));
    InMux I__452 (
            .O(N__2405),
            .I(N__2402));
    LocalMux I__451 (
            .O(N__2402),
            .I(N__2398));
    InMux I__450 (
            .O(N__2401),
            .I(N__2395));
    Odrv4 I__449 (
            .O(N__2398),
            .I(\Debounce_Sw1.un9_r_count_9 ));
    LocalMux I__448 (
            .O(N__2395),
            .I(\Debounce_Sw1.un9_r_count_9 ));
    InMux I__447 (
            .O(N__2390),
            .I(N__2385));
    InMux I__446 (
            .O(N__2389),
            .I(N__2382));
    InMux I__445 (
            .O(N__2388),
            .I(N__2379));
    LocalMux I__444 (
            .O(N__2385),
            .I(\Debounce_Sw1.r_CountZ0Z_12 ));
    LocalMux I__443 (
            .O(N__2382),
            .I(\Debounce_Sw1.r_CountZ0Z_12 ));
    LocalMux I__442 (
            .O(N__2379),
            .I(\Debounce_Sw1.r_CountZ0Z_12 ));
    InMux I__441 (
            .O(N__2372),
            .I(N__2367));
    InMux I__440 (
            .O(N__2371),
            .I(N__2364));
    InMux I__439 (
            .O(N__2370),
            .I(N__2361));
    LocalMux I__438 (
            .O(N__2367),
            .I(\Debounce_Sw1.r_CountZ0Z_14 ));
    LocalMux I__437 (
            .O(N__2364),
            .I(\Debounce_Sw1.r_CountZ0Z_14 ));
    LocalMux I__436 (
            .O(N__2361),
            .I(\Debounce_Sw1.r_CountZ0Z_14 ));
    CascadeMux I__435 (
            .O(N__2354),
            .I(N__2350));
    InMux I__434 (
            .O(N__2353),
            .I(N__2346));
    InMux I__433 (
            .O(N__2350),
            .I(N__2343));
    InMux I__432 (
            .O(N__2349),
            .I(N__2340));
    LocalMux I__431 (
            .O(N__2346),
            .I(\Debounce_Sw1.r_CountZ0Z_15 ));
    LocalMux I__430 (
            .O(N__2343),
            .I(\Debounce_Sw1.r_CountZ0Z_15 ));
    LocalMux I__429 (
            .O(N__2340),
            .I(\Debounce_Sw1.r_CountZ0Z_15 ));
    InMux I__428 (
            .O(N__2333),
            .I(N__2328));
    InMux I__427 (
            .O(N__2332),
            .I(N__2325));
    InMux I__426 (
            .O(N__2331),
            .I(N__2322));
    LocalMux I__425 (
            .O(N__2328),
            .I(\Debounce_Sw1.r_CountZ0Z_7 ));
    LocalMux I__424 (
            .O(N__2325),
            .I(\Debounce_Sw1.r_CountZ0Z_7 ));
    LocalMux I__423 (
            .O(N__2322),
            .I(\Debounce_Sw1.r_CountZ0Z_7 ));
    InMux I__422 (
            .O(N__2315),
            .I(N__2312));
    LocalMux I__421 (
            .O(N__2312),
            .I(N__2309));
    Odrv12 I__420 (
            .O(N__2309),
            .I(\Debounce_Sw1.un9_r_count_10 ));
    InMux I__419 (
            .O(N__2306),
            .I(N__2301));
    InMux I__418 (
            .O(N__2305),
            .I(N__2298));
    InMux I__417 (
            .O(N__2304),
            .I(N__2295));
    LocalMux I__416 (
            .O(N__2301),
            .I(\Debounce_Sw1.r_CountZ0Z_9 ));
    LocalMux I__415 (
            .O(N__2298),
            .I(\Debounce_Sw1.r_CountZ0Z_9 ));
    LocalMux I__414 (
            .O(N__2295),
            .I(\Debounce_Sw1.r_CountZ0Z_9 ));
    CascadeMux I__413 (
            .O(N__2288),
            .I(\Debounce_Sw1.un9_r_count_5_cascade_ ));
    InMux I__412 (
            .O(N__2285),
            .I(N__2280));
    InMux I__411 (
            .O(N__2284),
            .I(N__2277));
    InMux I__410 (
            .O(N__2283),
            .I(N__2274));
    LocalMux I__409 (
            .O(N__2280),
            .I(\Debounce_Sw1.r_CountZ0Z_10 ));
    LocalMux I__408 (
            .O(N__2277),
            .I(\Debounce_Sw1.r_CountZ0Z_10 ));
    LocalMux I__407 (
            .O(N__2274),
            .I(\Debounce_Sw1.r_CountZ0Z_10 ));
    InMux I__406 (
            .O(N__2267),
            .I(N__2264));
    LocalMux I__405 (
            .O(N__2264),
            .I(\Debounce_Sw1.un9_r_count_9_0 ));
    InMux I__404 (
            .O(N__2261),
            .I(N__2258));
    LocalMux I__403 (
            .O(N__2258),
            .I(N__2255));
    Span4Mux_h I__402 (
            .O(N__2255),
            .I(N__2251));
    InMux I__401 (
            .O(N__2254),
            .I(N__2248));
    Sp12to4 I__400 (
            .O(N__2251),
            .I(N__2243));
    LocalMux I__399 (
            .O(N__2248),
            .I(N__2243));
    Span12Mux_v I__398 (
            .O(N__2243),
            .I(N__2240));
    Odrv12 I__397 (
            .O(N__2240),
            .I(i_Switch_1_c));
    CascadeMux I__396 (
            .O(N__2237),
            .I(\Debounce_Sw1.un9_r_count_10_0_cascade_ ));
    InMux I__395 (
            .O(N__2234),
            .I(N__2229));
    InMux I__394 (
            .O(N__2233),
            .I(N__2226));
    InMux I__393 (
            .O(N__2232),
            .I(N__2223));
    LocalMux I__392 (
            .O(N__2229),
            .I(N__2220));
    LocalMux I__391 (
            .O(N__2226),
            .I(\Debounce_Sw1.r_CountZ0Z_16 ));
    LocalMux I__390 (
            .O(N__2223),
            .I(\Debounce_Sw1.r_CountZ0Z_16 ));
    Odrv4 I__389 (
            .O(N__2220),
            .I(\Debounce_Sw1.r_CountZ0Z_16 ));
    InMux I__388 (
            .O(N__2213),
            .I(N__2208));
    InMux I__387 (
            .O(N__2212),
            .I(N__2205));
    InMux I__386 (
            .O(N__2211),
            .I(N__2202));
    LocalMux I__385 (
            .O(N__2208),
            .I(\Debounce_Sw1.r_CountZ0Z_13 ));
    LocalMux I__384 (
            .O(N__2205),
            .I(\Debounce_Sw1.r_CountZ0Z_13 ));
    LocalMux I__383 (
            .O(N__2202),
            .I(\Debounce_Sw1.r_CountZ0Z_13 ));
    CascadeMux I__382 (
            .O(N__2195),
            .I(N__2191));
    CascadeMux I__381 (
            .O(N__2194),
            .I(N__2187));
    InMux I__380 (
            .O(N__2191),
            .I(N__2184));
    InMux I__379 (
            .O(N__2190),
            .I(N__2181));
    InMux I__378 (
            .O(N__2187),
            .I(N__2178));
    LocalMux I__377 (
            .O(N__2184),
            .I(N__2175));
    LocalMux I__376 (
            .O(N__2181),
            .I(\Debounce_Sw1.r_CountZ0Z_17 ));
    LocalMux I__375 (
            .O(N__2178),
            .I(\Debounce_Sw1.r_CountZ0Z_17 ));
    Odrv4 I__374 (
            .O(N__2175),
            .I(\Debounce_Sw1.r_CountZ0Z_17 ));
    CascadeMux I__373 (
            .O(N__2168),
            .I(N__2163));
    InMux I__372 (
            .O(N__2167),
            .I(N__2160));
    InMux I__371 (
            .O(N__2166),
            .I(N__2157));
    InMux I__370 (
            .O(N__2163),
            .I(N__2154));
    LocalMux I__369 (
            .O(N__2160),
            .I(\Debounce_Sw1.r_CountZ0Z_11 ));
    LocalMux I__368 (
            .O(N__2157),
            .I(\Debounce_Sw1.r_CountZ0Z_11 ));
    LocalMux I__367 (
            .O(N__2154),
            .I(\Debounce_Sw1.r_CountZ0Z_11 ));
    InMux I__366 (
            .O(N__2147),
            .I(N__2144));
    LocalMux I__365 (
            .O(N__2144),
            .I(\Debounce_Sw1.un9_r_count_6 ));
    InMux I__364 (
            .O(N__2141),
            .I(N__2138));
    LocalMux I__363 (
            .O(N__2138),
            .I(N__2135));
    Odrv4 I__362 (
            .O(N__2135),
            .I(\Count_And_Toggle.r_Counter_RNO_0Z0Z_9 ));
    CascadeMux I__361 (
            .O(N__2132),
            .I(N__2128));
    InMux I__360 (
            .O(N__2131),
            .I(N__2125));
    InMux I__359 (
            .O(N__2128),
            .I(N__2122));
    LocalMux I__358 (
            .O(N__2125),
            .I(N__2119));
    LocalMux I__357 (
            .O(N__2122),
            .I(\Count_And_Toggle.r_CounterZ0Z_9 ));
    Odrv4 I__356 (
            .O(N__2119),
            .I(\Count_And_Toggle.r_CounterZ0Z_9 ));
    CascadeMux I__355 (
            .O(N__2114),
            .I(N__2111));
    InMux I__354 (
            .O(N__2111),
            .I(N__2106));
    CascadeMux I__353 (
            .O(N__2110),
            .I(N__2101));
    CascadeMux I__352 (
            .O(N__2109),
            .I(N__2097));
    LocalMux I__351 (
            .O(N__2106),
            .I(N__2094));
    InMux I__350 (
            .O(N__2105),
            .I(N__2091));
    CascadeMux I__349 (
            .O(N__2104),
            .I(N__2087));
    InMux I__348 (
            .O(N__2101),
            .I(N__2078));
    InMux I__347 (
            .O(N__2100),
            .I(N__2078));
    InMux I__346 (
            .O(N__2097),
            .I(N__2078));
    Span4Mux_v I__345 (
            .O(N__2094),
            .I(N__2073));
    LocalMux I__344 (
            .O(N__2091),
            .I(N__2073));
    InMux I__343 (
            .O(N__2090),
            .I(N__2070));
    InMux I__342 (
            .O(N__2087),
            .I(N__2065));
    InMux I__341 (
            .O(N__2086),
            .I(N__2065));
    InMux I__340 (
            .O(N__2085),
            .I(N__2062));
    LocalMux I__339 (
            .O(N__2078),
            .I(\Count_And_Toggle.un4_i_enable_16 ));
    Odrv4 I__338 (
            .O(N__2073),
            .I(\Count_And_Toggle.un4_i_enable_16 ));
    LocalMux I__337 (
            .O(N__2070),
            .I(\Count_And_Toggle.un4_i_enable_16 ));
    LocalMux I__336 (
            .O(N__2065),
            .I(\Count_And_Toggle.un4_i_enable_16 ));
    LocalMux I__335 (
            .O(N__2062),
            .I(\Count_And_Toggle.un4_i_enable_16 ));
    CascadeMux I__334 (
            .O(N__2051),
            .I(N__2045));
    InMux I__333 (
            .O(N__2050),
            .I(N__2038));
    InMux I__332 (
            .O(N__2049),
            .I(N__2035));
    InMux I__331 (
            .O(N__2048),
            .I(N__2028));
    InMux I__330 (
            .O(N__2045),
            .I(N__2028));
    InMux I__329 (
            .O(N__2044),
            .I(N__2028));
    InMux I__328 (
            .O(N__2043),
            .I(N__2025));
    InMux I__327 (
            .O(N__2042),
            .I(N__2020));
    InMux I__326 (
            .O(N__2041),
            .I(N__2020));
    LocalMux I__325 (
            .O(N__2038),
            .I(\Count_And_Toggle.un4_i_enable_15 ));
    LocalMux I__324 (
            .O(N__2035),
            .I(\Count_And_Toggle.un4_i_enable_15 ));
    LocalMux I__323 (
            .O(N__2028),
            .I(\Count_And_Toggle.un4_i_enable_15 ));
    LocalMux I__322 (
            .O(N__2025),
            .I(\Count_And_Toggle.un4_i_enable_15 ));
    LocalMux I__321 (
            .O(N__2020),
            .I(\Count_And_Toggle.un4_i_enable_15 ));
    InMux I__320 (
            .O(N__2009),
            .I(N__2006));
    LocalMux I__319 (
            .O(N__2006),
            .I(\Count_And_Toggle.r_Counter_RNO_0Z0Z_11 ));
    InMux I__318 (
            .O(N__2003),
            .I(N__1999));
    InMux I__317 (
            .O(N__2002),
            .I(N__1996));
    LocalMux I__316 (
            .O(N__1999),
            .I(\Count_And_Toggle.r_CounterZ0Z_3 ));
    LocalMux I__315 (
            .O(N__1996),
            .I(\Count_And_Toggle.r_CounterZ0Z_3 ));
    InMux I__314 (
            .O(N__1991),
            .I(N__1987));
    InMux I__313 (
            .O(N__1990),
            .I(N__1984));
    LocalMux I__312 (
            .O(N__1987),
            .I(\Count_And_Toggle.r_CounterZ0Z_2 ));
    LocalMux I__311 (
            .O(N__1984),
            .I(\Count_And_Toggle.r_CounterZ0Z_2 ));
    InMux I__310 (
            .O(N__1979),
            .I(N__1972));
    InMux I__309 (
            .O(N__1978),
            .I(N__1972));
    InMux I__308 (
            .O(N__1977),
            .I(N__1969));
    LocalMux I__307 (
            .O(N__1972),
            .I(\Count_And_Toggle.r_CounterZ0Z_1 ));
    LocalMux I__306 (
            .O(N__1969),
            .I(\Count_And_Toggle.r_CounterZ0Z_1 ));
    InMux I__305 (
            .O(N__1964),
            .I(N__1961));
    LocalMux I__304 (
            .O(N__1961),
            .I(N__1958));
    Odrv4 I__303 (
            .O(N__1958),
            .I(\Count_And_Toggle.r_Counter_RNO_0Z0Z_6 ));
    CascadeMux I__302 (
            .O(N__1955),
            .I(N__1952));
    InMux I__301 (
            .O(N__1952),
            .I(N__1948));
    InMux I__300 (
            .O(N__1951),
            .I(N__1945));
    LocalMux I__299 (
            .O(N__1948),
            .I(\Count_And_Toggle.r_CounterZ0Z_6 ));
    LocalMux I__298 (
            .O(N__1945),
            .I(\Count_And_Toggle.r_CounterZ0Z_6 ));
    InMux I__297 (
            .O(N__1940),
            .I(N__1937));
    LocalMux I__296 (
            .O(N__1937),
            .I(\Count_And_Toggle.r_Counter_RNO_0Z0Z_19 ));
    CascadeMux I__295 (
            .O(N__1934),
            .I(N__1930));
    CascadeMux I__294 (
            .O(N__1933),
            .I(N__1927));
    InMux I__293 (
            .O(N__1930),
            .I(N__1924));
    InMux I__292 (
            .O(N__1927),
            .I(N__1921));
    LocalMux I__291 (
            .O(N__1924),
            .I(\Count_And_Toggle.r_CounterZ0Z_19 ));
    LocalMux I__290 (
            .O(N__1921),
            .I(\Count_And_Toggle.r_CounterZ0Z_19 ));
    InMux I__289 (
            .O(N__1916),
            .I(N__1912));
    InMux I__288 (
            .O(N__1915),
            .I(N__1909));
    LocalMux I__287 (
            .O(N__1912),
            .I(\Count_And_Toggle.r_CounterZ0Z_11 ));
    LocalMux I__286 (
            .O(N__1909),
            .I(\Count_And_Toggle.r_CounterZ0Z_11 ));
    CascadeMux I__285 (
            .O(N__1904),
            .I(\Count_And_Toggle.un4_i_enable_15_cascade_ ));
    InMux I__284 (
            .O(N__1901),
            .I(N__1898));
    LocalMux I__283 (
            .O(N__1898),
            .I(\Count_And_Toggle.r_Counter_RNO_0Z0Z_18 ));
    InMux I__282 (
            .O(N__1895),
            .I(N__1891));
    InMux I__281 (
            .O(N__1894),
            .I(N__1888));
    LocalMux I__280 (
            .O(N__1891),
            .I(\Count_And_Toggle.r_CounterZ0Z_18 ));
    LocalMux I__279 (
            .O(N__1888),
            .I(\Count_And_Toggle.r_CounterZ0Z_18 ));
    InMux I__278 (
            .O(N__1883),
            .I(N__1879));
    InMux I__277 (
            .O(N__1882),
            .I(N__1876));
    LocalMux I__276 (
            .O(N__1879),
            .I(\Count_And_Toggle.r_CounterZ0Z_15 ));
    LocalMux I__275 (
            .O(N__1876),
            .I(\Count_And_Toggle.r_CounterZ0Z_15 ));
    InMux I__274 (
            .O(N__1871),
            .I(N__1867));
    InMux I__273 (
            .O(N__1870),
            .I(N__1864));
    LocalMux I__272 (
            .O(N__1867),
            .I(\Count_And_Toggle.r_CounterZ0Z_16 ));
    LocalMux I__271 (
            .O(N__1864),
            .I(\Count_And_Toggle.r_CounterZ0Z_16 ));
    CascadeMux I__270 (
            .O(N__1859),
            .I(N__1853));
    InMux I__269 (
            .O(N__1858),
            .I(N__1848));
    InMux I__268 (
            .O(N__1857),
            .I(N__1848));
    InMux I__267 (
            .O(N__1856),
            .I(N__1845));
    InMux I__266 (
            .O(N__1853),
            .I(N__1842));
    LocalMux I__265 (
            .O(N__1848),
            .I(\Count_And_Toggle.r_CounterZ0Z_0 ));
    LocalMux I__264 (
            .O(N__1845),
            .I(\Count_And_Toggle.r_CounterZ0Z_0 ));
    LocalMux I__263 (
            .O(N__1842),
            .I(\Count_And_Toggle.r_CounterZ0Z_0 ));
    InMux I__262 (
            .O(N__1835),
            .I(N__1832));
    LocalMux I__261 (
            .O(N__1832),
            .I(\Count_And_Toggle.un4_i_enable_14 ));
    InMux I__260 (
            .O(N__1829),
            .I(N__1826));
    LocalMux I__259 (
            .O(N__1826),
            .I(\Count_And_Toggle.un4_i_enable_12 ));
    CascadeMux I__258 (
            .O(N__1823),
            .I(\Count_And_Toggle.un4_i_enable_11_cascade_ ));
    InMux I__257 (
            .O(N__1820),
            .I(N__1817));
    LocalMux I__256 (
            .O(N__1817),
            .I(\Count_And_Toggle.un4_i_enable_13 ));
    InMux I__255 (
            .O(N__1814),
            .I(\Debounce_Sw1.un2_r_count_cry_13 ));
    InMux I__254 (
            .O(N__1811),
            .I(\Debounce_Sw1.un2_r_count_cry_14 ));
    InMux I__253 (
            .O(N__1808),
            .I(\Debounce_Sw1.un2_r_count_cry_15 ));
    InMux I__252 (
            .O(N__1805),
            .I(bfn_5_7_0_));
    SRMux I__251 (
            .O(N__1802),
            .I(N__1790));
    SRMux I__250 (
            .O(N__1801),
            .I(N__1790));
    SRMux I__249 (
            .O(N__1800),
            .I(N__1790));
    SRMux I__248 (
            .O(N__1799),
            .I(N__1790));
    GlobalMux I__247 (
            .O(N__1790),
            .I(N__1787));
    gio2CtrlBuf I__246 (
            .O(N__1787),
            .I(\Debounce_Sw1.r_count15_i_g ));
    InMux I__245 (
            .O(N__1784),
            .I(N__1781));
    LocalMux I__244 (
            .O(N__1781),
            .I(N__1777));
    InMux I__243 (
            .O(N__1780),
            .I(N__1774));
    Odrv4 I__242 (
            .O(N__1777),
            .I(\Count_And_Toggle.r_CounterZ0Z_12 ));
    LocalMux I__241 (
            .O(N__1774),
            .I(\Count_And_Toggle.r_CounterZ0Z_12 ));
    InMux I__240 (
            .O(N__1769),
            .I(N__1765));
    InMux I__239 (
            .O(N__1768),
            .I(N__1762));
    LocalMux I__238 (
            .O(N__1765),
            .I(\Count_And_Toggle.r_CounterZ0Z_10 ));
    LocalMux I__237 (
            .O(N__1762),
            .I(\Count_And_Toggle.r_CounterZ0Z_10 ));
    CascadeMux I__236 (
            .O(N__1757),
            .I(N__1754));
    InMux I__235 (
            .O(N__1754),
            .I(N__1750));
    InMux I__234 (
            .O(N__1753),
            .I(N__1747));
    LocalMux I__233 (
            .O(N__1750),
            .I(\Count_And_Toggle.r_CounterZ0Z_13 ));
    LocalMux I__232 (
            .O(N__1747),
            .I(\Count_And_Toggle.r_CounterZ0Z_13 ));
    InMux I__231 (
            .O(N__1742),
            .I(N__1738));
    InMux I__230 (
            .O(N__1741),
            .I(N__1735));
    LocalMux I__229 (
            .O(N__1738),
            .I(\Count_And_Toggle.r_CounterZ0Z_7 ));
    LocalMux I__228 (
            .O(N__1735),
            .I(\Count_And_Toggle.r_CounterZ0Z_7 ));
    InMux I__227 (
            .O(N__1730),
            .I(N__1727));
    LocalMux I__226 (
            .O(N__1727),
            .I(\Count_And_Toggle.r_Counter_RNO_0Z0Z_8 ));
    CascadeMux I__225 (
            .O(N__1724),
            .I(N__1720));
    InMux I__224 (
            .O(N__1723),
            .I(N__1717));
    InMux I__223 (
            .O(N__1720),
            .I(N__1714));
    LocalMux I__222 (
            .O(N__1717),
            .I(\Count_And_Toggle.r_CounterZ0Z_8 ));
    LocalMux I__221 (
            .O(N__1714),
            .I(\Count_And_Toggle.r_CounterZ0Z_8 ));
    InMux I__220 (
            .O(N__1709),
            .I(N__1705));
    InMux I__219 (
            .O(N__1708),
            .I(N__1702));
    LocalMux I__218 (
            .O(N__1705),
            .I(\Count_And_Toggle.r_CounterZ0Z_5 ));
    LocalMux I__217 (
            .O(N__1702),
            .I(\Count_And_Toggle.r_CounterZ0Z_5 ));
    InMux I__216 (
            .O(N__1697),
            .I(N__1693));
    InMux I__215 (
            .O(N__1696),
            .I(N__1690));
    LocalMux I__214 (
            .O(N__1693),
            .I(\Count_And_Toggle.r_CounterZ0Z_4 ));
    LocalMux I__213 (
            .O(N__1690),
            .I(\Count_And_Toggle.r_CounterZ0Z_4 ));
    InMux I__212 (
            .O(N__1685),
            .I(N__1681));
    InMux I__211 (
            .O(N__1684),
            .I(N__1678));
    LocalMux I__210 (
            .O(N__1681),
            .I(\Debounce_Sw1.r_CountZ0Z_5 ));
    LocalMux I__209 (
            .O(N__1678),
            .I(\Debounce_Sw1.r_CountZ0Z_5 ));
    InMux I__208 (
            .O(N__1673),
            .I(\Debounce_Sw1.un2_r_count_cry_4 ));
    InMux I__207 (
            .O(N__1670),
            .I(\Debounce_Sw1.un2_r_count_cry_5 ));
    InMux I__206 (
            .O(N__1667),
            .I(\Debounce_Sw1.un2_r_count_cry_6 ));
    InMux I__205 (
            .O(N__1664),
            .I(\Debounce_Sw1.un2_r_count_cry_7 ));
    InMux I__204 (
            .O(N__1661),
            .I(bfn_5_6_0_));
    InMux I__203 (
            .O(N__1658),
            .I(\Debounce_Sw1.un2_r_count_cry_9 ));
    InMux I__202 (
            .O(N__1655),
            .I(\Debounce_Sw1.un2_r_count_cry_10 ));
    InMux I__201 (
            .O(N__1652),
            .I(\Debounce_Sw1.un2_r_count_cry_11 ));
    InMux I__200 (
            .O(N__1649),
            .I(\Debounce_Sw1.un2_r_count_cry_12 ));
    InMux I__199 (
            .O(N__1646),
            .I(\Count_And_Toggle.un2_r_counter_cry_19 ));
    InMux I__198 (
            .O(N__1643),
            .I(\Count_And_Toggle.un2_r_counter_cry_20 ));
    InMux I__197 (
            .O(N__1640),
            .I(\Count_And_Toggle.un2_r_counter_cry_21 ));
    CascadeMux I__196 (
            .O(N__1637),
            .I(\Count_And_Toggle.r_Counter_RNO_0Z0Z_22_cascade_ ));
    InMux I__195 (
            .O(N__1634),
            .I(N__1628));
    InMux I__194 (
            .O(N__1633),
            .I(N__1628));
    LocalMux I__193 (
            .O(N__1628),
            .I(\Count_And_Toggle.r_CounterZ0Z_17 ));
    InMux I__192 (
            .O(N__1625),
            .I(N__1619));
    InMux I__191 (
            .O(N__1624),
            .I(N__1619));
    LocalMux I__190 (
            .O(N__1619),
            .I(\Count_And_Toggle.r_CounterZ0Z_22 ));
    CascadeMux I__189 (
            .O(N__1616),
            .I(N__1613));
    InMux I__188 (
            .O(N__1613),
            .I(N__1607));
    InMux I__187 (
            .O(N__1612),
            .I(N__1607));
    LocalMux I__186 (
            .O(N__1607),
            .I(\Count_And_Toggle.r_CounterZ0Z_21 ));
    InMux I__185 (
            .O(N__1604),
            .I(N__1598));
    InMux I__184 (
            .O(N__1603),
            .I(N__1598));
    LocalMux I__183 (
            .O(N__1598),
            .I(\Count_And_Toggle.r_CounterZ0Z_20 ));
    InMux I__182 (
            .O(N__1595),
            .I(N__1589));
    InMux I__181 (
            .O(N__1594),
            .I(N__1582));
    InMux I__180 (
            .O(N__1593),
            .I(N__1582));
    InMux I__179 (
            .O(N__1592),
            .I(N__1582));
    LocalMux I__178 (
            .O(N__1589),
            .I(\Debounce_Sw1.r_CountZ0Z_0 ));
    LocalMux I__177 (
            .O(N__1582),
            .I(\Debounce_Sw1.r_CountZ0Z_0 ));
    CascadeMux I__176 (
            .O(N__1577),
            .I(N__1573));
    CascadeMux I__175 (
            .O(N__1576),
            .I(N__1570));
    InMux I__174 (
            .O(N__1573),
            .I(N__1566));
    InMux I__173 (
            .O(N__1570),
            .I(N__1561));
    InMux I__172 (
            .O(N__1569),
            .I(N__1561));
    LocalMux I__171 (
            .O(N__1566),
            .I(\Debounce_Sw1.r_CountZ0Z_1 ));
    LocalMux I__170 (
            .O(N__1561),
            .I(\Debounce_Sw1.r_CountZ0Z_1 ));
    InMux I__169 (
            .O(N__1556),
            .I(N__1552));
    InMux I__168 (
            .O(N__1555),
            .I(N__1549));
    LocalMux I__167 (
            .O(N__1552),
            .I(\Debounce_Sw1.r_CountZ0Z_2 ));
    LocalMux I__166 (
            .O(N__1549),
            .I(\Debounce_Sw1.r_CountZ0Z_2 ));
    InMux I__165 (
            .O(N__1544),
            .I(\Debounce_Sw1.un2_r_count_cry_1 ));
    CascadeMux I__164 (
            .O(N__1541),
            .I(N__1537));
    InMux I__163 (
            .O(N__1540),
            .I(N__1534));
    InMux I__162 (
            .O(N__1537),
            .I(N__1531));
    LocalMux I__161 (
            .O(N__1534),
            .I(\Debounce_Sw1.r_CountZ0Z_3 ));
    LocalMux I__160 (
            .O(N__1531),
            .I(\Debounce_Sw1.r_CountZ0Z_3 ));
    InMux I__159 (
            .O(N__1526),
            .I(\Debounce_Sw1.un2_r_count_cry_2 ));
    InMux I__158 (
            .O(N__1523),
            .I(N__1519));
    InMux I__157 (
            .O(N__1522),
            .I(N__1516));
    LocalMux I__156 (
            .O(N__1519),
            .I(\Debounce_Sw1.r_CountZ0Z_4 ));
    LocalMux I__155 (
            .O(N__1516),
            .I(\Debounce_Sw1.r_CountZ0Z_4 ));
    InMux I__154 (
            .O(N__1511),
            .I(\Debounce_Sw1.un2_r_count_cry_3 ));
    InMux I__153 (
            .O(N__1508),
            .I(\Count_And_Toggle.un2_r_counter_cry_10 ));
    InMux I__152 (
            .O(N__1505),
            .I(\Count_And_Toggle.un2_r_counter_cry_11 ));
    InMux I__151 (
            .O(N__1502),
            .I(\Count_And_Toggle.un2_r_counter_cry_12 ));
    InMux I__150 (
            .O(N__1499),
            .I(\Count_And_Toggle.un2_r_counter_cry_13 ));
    InMux I__149 (
            .O(N__1496),
            .I(\Count_And_Toggle.un2_r_counter_cry_14 ));
    InMux I__148 (
            .O(N__1493),
            .I(\Count_And_Toggle.un2_r_counter_cry_15 ));
    InMux I__147 (
            .O(N__1490),
            .I(bfn_4_9_0_));
    InMux I__146 (
            .O(N__1487),
            .I(\Count_And_Toggle.un2_r_counter_cry_17 ));
    InMux I__145 (
            .O(N__1484),
            .I(\Count_And_Toggle.un2_r_counter_cry_18 ));
    InMux I__144 (
            .O(N__1481),
            .I(\Count_And_Toggle.un2_r_counter_cry_1 ));
    InMux I__143 (
            .O(N__1478),
            .I(\Count_And_Toggle.un2_r_counter_cry_2 ));
    InMux I__142 (
            .O(N__1475),
            .I(\Count_And_Toggle.un2_r_counter_cry_3 ));
    InMux I__141 (
            .O(N__1472),
            .I(\Count_And_Toggle.un2_r_counter_cry_4 ));
    InMux I__140 (
            .O(N__1469),
            .I(\Count_And_Toggle.un2_r_counter_cry_5 ));
    InMux I__139 (
            .O(N__1466),
            .I(\Count_And_Toggle.un2_r_counter_cry_6 ));
    InMux I__138 (
            .O(N__1463),
            .I(\Count_And_Toggle.un2_r_counter_cry_7 ));
    InMux I__137 (
            .O(N__1460),
            .I(bfn_4_8_0_));
    InMux I__136 (
            .O(N__1457),
            .I(\Count_And_Toggle.un2_r_counter_cry_9 ));
    CascadeMux I__135 (
            .O(N__1454),
            .I(\Debounce_Sw1.un9_r_count_10_cascade_ ));
    CascadeMux I__134 (
            .O(N__1451),
            .I(\Debounce_Sw1.un1_r_Count_1lt11_0_cascade_ ));
    InMux I__133 (
            .O(N__1448),
            .I(N__1445));
    LocalMux I__132 (
            .O(N__1445),
            .I(\Debounce_Sw1.un1_r_Count_1lto11_1 ));
    CascadeMux I__131 (
            .O(N__1442),
            .I(\Debounce_Sw1.un1_r_Count_1lt17_cascade_ ));
    InMux I__130 (
            .O(N__1439),
            .I(N__1436));
    LocalMux I__129 (
            .O(N__1436),
            .I(\Debounce_Sw1.un1_r_Count_1lto17_2 ));
    IoInMux I__128 (
            .O(N__1433),
            .I(N__1430));
    LocalMux I__127 (
            .O(N__1430),
            .I(N__1427));
    Span4Mux_s3_h I__126 (
            .O(N__1427),
            .I(N__1424));
    Odrv4 I__125 (
            .O(N__1424),
            .I(\Debounce_Sw1.r_count15_i ));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\Debounce_Sw2.un2_r_count_cry_8 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(\Debounce_Sw2.un2_r_count_cry_16 ),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_5_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_5_0_));
    defparam IN_MUX_bfv_5_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_6_0_ (
            .carryinitin(\Debounce_Sw1.un2_r_count_cry_8 ),
            .carryinitout(bfn_5_6_0_));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(\Debounce_Sw1.un2_r_count_cry_16 ),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_4_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_7_0_));
    defparam IN_MUX_bfv_4_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_8_0_ (
            .carryinitin(\Count_And_Toggle.un2_r_counter_cry_8 ),
            .carryinitout(bfn_4_8_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(\Count_And_Toggle.un2_r_counter_cry_16 ),
            .carryinitout(bfn_4_9_0_));
    ICE_GB \Debounce_Sw2.r_State_e_0_RNIK82U4_0  (
            .USERSIGNALTOGLOBALBUFFER(N__2495),
            .GLOBALBUFFEROUTPUT(\Debounce_Sw2.N_9_g ));
    ICE_GB \Debounce_Sw1.r_State_RNIDSE73_0  (
            .USERSIGNALTOGLOBALBUFFER(N__1433),
            .GLOBALBUFFEROUTPUT(\Debounce_Sw1.r_count15_i_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \Debounce_Sw1.r_Count_RNI720A_4_LC_4_5_3 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_Count_RNI720A_4_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw1.r_Count_RNI720A_4_LC_4_5_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Debounce_Sw1.r_Count_RNI720A_4_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(N__1522),
            .in2(_gnd_net_),
            .in3(N__1684),
            .lcout(\Debounce_Sw1.un9_r_count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.r_Count_RNIGFOJ_10_LC_4_5_5 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_Count_RNIGFOJ_10_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw1.r_Count_RNIGFOJ_10_LC_4_5_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Debounce_Sw1.r_Count_RNIGFOJ_10_LC_4_5_5  (
            .in0(N__2283),
            .in1(N__2304),
            .in2(N__2168),
            .in3(N__2442),
            .lcout(\Debounce_Sw1.un1_r_Count_1lto11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.r_Count_RNIMUGJ_17_LC_4_5_6 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_Count_RNIMUGJ_17_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw1.r_Count_RNIMUGJ_17_LC_4_5_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_Sw1.r_Count_RNIMUGJ_17_LC_4_5_6  (
            .in0(N__2234),
            .in1(N__2349),
            .in2(N__2195),
            .in3(N__2370),
            .lcout(\Debounce_Sw1.un1_r_Count_1lto17_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.r_Count_1_LC_4_6_2 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_Count_1_LC_4_6_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_1_LC_4_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Debounce_Sw1.r_Count_1_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1576),
            .in3(N__1593),
            .lcout(\Debounce_Sw1.r_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3075),
            .ce(),
            .sr(N__1799));
    defparam \Debounce_Sw1.r_Count_RNI2OVJ_1_LC_4_6_3 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_Count_RNI2OVJ_1_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw1.r_Count_RNI2OVJ_1_LC_4_6_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_Sw1.r_Count_RNI2OVJ_1_LC_4_6_3  (
            .in0(N__1592),
            .in1(N__1569),
            .in2(N__1541),
            .in3(N__1555),
            .lcout(\Debounce_Sw1.un9_r_count_10 ),
            .ltout(\Debounce_Sw1.un9_r_count_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.r_Count_RNIK0081_6_LC_4_6_4 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_Count_RNIK0081_6_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw1.r_Count_RNIK0081_6_LC_4_6_4 .LUT_INIT=16'b1010100010101010;
    LogicCell40 \Debounce_Sw1.r_Count_RNIK0081_6_LC_4_6_4  (
            .in0(N__2331),
            .in1(N__2421),
            .in2(N__1454),
            .in3(N__2401),
            .lcout(),
            .ltout(\Debounce_Sw1.un1_r_Count_1lt11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.r_Count_RNI9PG52_12_LC_4_6_5 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_Count_RNI9PG52_12_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw1.r_Count_RNI9PG52_12_LC_4_6_5 .LUT_INIT=16'b0001010100010001;
    LogicCell40 \Debounce_Sw1.r_Count_RNI9PG52_12_LC_4_6_5  (
            .in0(N__2211),
            .in1(N__2388),
            .in2(N__1451),
            .in3(N__1448),
            .lcout(),
            .ltout(\Debounce_Sw1.un1_r_Count_1lt17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.r_State_RNIDSE73_LC_4_6_6 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_State_RNIDSE73_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw1.r_State_RNIDSE73_LC_4_6_6 .LUT_INIT=16'b1001111110011001;
    LogicCell40 \Debounce_Sw1.r_State_RNIDSE73_LC_4_6_6  (
            .in0(N__2261),
            .in1(N__2974),
            .in2(N__1442),
            .in3(N__1439),
            .lcout(\Debounce_Sw1.r_count15_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.r_Count_0_LC_4_6_7 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_Count_0_LC_4_6_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_0_LC_4_6_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \Debounce_Sw1.r_Count_0_LC_4_6_7  (
            .in0(N__1594),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Debounce_Sw1.r_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3075),
            .ce(),
            .sr(N__1799));
    defparam \Count_And_Toggle.un2_r_counter_cry_1_c_LC_4_7_0 .C_ON=1'b1;
    defparam \Count_And_Toggle.un2_r_counter_cry_1_c_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.un2_r_counter_cry_1_c_LC_4_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Count_And_Toggle.un2_r_counter_cry_1_c_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(N__1977),
            .in2(N__1859),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_7_0_),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_2_LC_4_7_1 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_2_LC_4_7_1 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_2_LC_4_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_2_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(N__1990),
            .in2(_gnd_net_),
            .in3(N__1481),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_2 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_1 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_2 ),
            .clk(N__3072),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_3_LC_4_7_2 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_3_LC_4_7_2 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_3_LC_4_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_3_LC_4_7_2  (
            .in0(_gnd_net_),
            .in1(N__2002),
            .in2(_gnd_net_),
            .in3(N__1478),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_3 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_2 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_3 ),
            .clk(N__3072),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_4_LC_4_7_3 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_4_LC_4_7_3 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_4_LC_4_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_4_LC_4_7_3  (
            .in0(_gnd_net_),
            .in1(N__1696),
            .in2(_gnd_net_),
            .in3(N__1475),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_4 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_3 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_4 ),
            .clk(N__3072),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_5_LC_4_7_4 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_5_LC_4_7_4 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_5_LC_4_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_5_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(N__1708),
            .in2(_gnd_net_),
            .in3(N__1472),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_5 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_4 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_5 ),
            .clk(N__3072),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNO_0_6_LC_4_7_5 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_RNO_0_6_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNO_0_6_LC_4_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_RNO_0_6_LC_4_7_5  (
            .in0(_gnd_net_),
            .in1(N__1951),
            .in2(_gnd_net_),
            .in3(N__1469),
            .lcout(\Count_And_Toggle.r_Counter_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_5 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_7_LC_4_7_6 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_7_LC_4_7_6 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_7_LC_4_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_7_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(N__1741),
            .in2(_gnd_net_),
            .in3(N__1466),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_7 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_6 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_7 ),
            .clk(N__3072),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNO_0_8_LC_4_7_7 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_RNO_0_8_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNO_0_8_LC_4_7_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Count_And_Toggle.r_Counter_RNO_0_8_LC_4_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1724),
            .in3(N__1463),
            .lcout(\Count_And_Toggle.r_Counter_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_7 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNO_0_9_LC_4_8_0 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_RNO_0_9_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNO_0_9_LC_4_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_RNO_0_9_LC_4_8_0  (
            .in0(_gnd_net_),
            .in1(N__2131),
            .in2(_gnd_net_),
            .in3(N__1460),
            .lcout(\Count_And_Toggle.r_Counter_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_4_8_0_),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_10_LC_4_8_1 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_10_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_10_LC_4_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_10_LC_4_8_1  (
            .in0(_gnd_net_),
            .in1(N__1768),
            .in2(_gnd_net_),
            .in3(N__1457),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_10 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_9 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_10 ),
            .clk(N__3070),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNO_0_11_LC_4_8_2 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_RNO_0_11_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNO_0_11_LC_4_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_RNO_0_11_LC_4_8_2  (
            .in0(_gnd_net_),
            .in1(N__1915),
            .in2(_gnd_net_),
            .in3(N__1508),
            .lcout(\Count_And_Toggle.r_Counter_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_10 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_12_LC_4_8_3 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_12_LC_4_8_3 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_12_LC_4_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_12_LC_4_8_3  (
            .in0(_gnd_net_),
            .in1(N__1780),
            .in2(_gnd_net_),
            .in3(N__1505),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_12 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_11 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_12 ),
            .clk(N__3070),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_13_LC_4_8_4 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_13_LC_4_8_4 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_13_LC_4_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_13_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(N__1753),
            .in2(_gnd_net_),
            .in3(N__1502),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_13 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_12 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_13 ),
            .clk(N__3070),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNO_0_14_LC_4_8_5 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_RNO_0_14_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNO_0_14_LC_4_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_RNO_0_14_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(N__2455),
            .in2(_gnd_net_),
            .in3(N__1499),
            .lcout(\Count_And_Toggle.r_Counter_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_13 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_15_LC_4_8_6 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_15_LC_4_8_6 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_15_LC_4_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_15_LC_4_8_6  (
            .in0(_gnd_net_),
            .in1(N__1882),
            .in2(_gnd_net_),
            .in3(N__1496),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_15 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_14 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_15 ),
            .clk(N__3070),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_16_LC_4_8_7 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_16_LC_4_8_7 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_16_LC_4_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_16_LC_4_8_7  (
            .in0(_gnd_net_),
            .in1(N__1870),
            .in2(_gnd_net_),
            .in3(N__1493),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_16 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_15 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_16 ),
            .clk(N__3070),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_17_LC_4_9_0 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_17_LC_4_9_0 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_17_LC_4_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_17_LC_4_9_0  (
            .in0(_gnd_net_),
            .in1(N__1633),
            .in2(_gnd_net_),
            .in3(N__1490),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_17 ),
            .clk(N__3073),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNO_0_18_LC_4_9_1 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_RNO_0_18_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNO_0_18_LC_4_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_RNO_0_18_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(N__1894),
            .in2(_gnd_net_),
            .in3(N__1487),
            .lcout(\Count_And_Toggle.r_Counter_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_17 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNO_0_19_LC_4_9_2 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_RNO_0_19_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNO_0_19_LC_4_9_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Count_And_Toggle.r_Counter_RNO_0_19_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1933),
            .in3(N__1484),
            .lcout(\Count_And_Toggle.r_Counter_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_18 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_20_LC_4_9_3 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_20_LC_4_9_3 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_20_LC_4_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_20_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__1603),
            .in2(_gnd_net_),
            .in3(N__1646),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_20 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_19 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_20 ),
            .clk(N__3073),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_21_LC_4_9_4 .C_ON=1'b1;
    defparam \Count_And_Toggle.r_Counter_21_LC_4_9_4 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_21_LC_4_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Count_And_Toggle.r_Counter_21_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(N__1612),
            .in2(_gnd_net_),
            .in3(N__1643),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_21 ),
            .ltout(),
            .carryin(\Count_And_Toggle.un2_r_counter_cry_20 ),
            .carryout(\Count_And_Toggle.un2_r_counter_cry_21 ),
            .clk(N__3073),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNO_0_22_LC_4_9_5 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_RNO_0_22_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNO_0_22_LC_4_9_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Count_And_Toggle.r_Counter_RNO_0_22_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(N__1625),
            .in2(_gnd_net_),
            .in3(N__1640),
            .lcout(),
            .ltout(\Count_And_Toggle.r_Counter_RNO_0Z0Z_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_22_LC_4_9_6 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_22_LC_4_9_6 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_22_LC_4_9_6 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \Count_And_Toggle.r_Counter_22_LC_4_9_6  (
            .in0(N__2085),
            .in1(N__2049),
            .in2(N__1637),
            .in3(N__2572),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3073),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNITEQL1_22_LC_4_9_7 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_RNITEQL1_22_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNITEQL1_22_LC_4_9_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Count_And_Toggle.r_Counter_RNITEQL1_22_LC_4_9_7  (
            .in0(N__1634),
            .in1(N__1624),
            .in2(N__1616),
            .in3(N__1604),
            .lcout(\Count_And_Toggle.un4_i_enable_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.un2_r_count_cry_1_c_LC_5_5_0 .C_ON=1'b1;
    defparam \Debounce_Sw1.un2_r_count_cry_1_c_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw1.un2_r_count_cry_1_c_LC_5_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Debounce_Sw1.un2_r_count_cry_1_c_LC_5_5_0  (
            .in0(_gnd_net_),
            .in1(N__1595),
            .in2(N__1577),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_5_0_),
            .carryout(\Debounce_Sw1.un2_r_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.r_Count_2_LC_5_5_1 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_2_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_2_LC_5_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_2_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(N__1556),
            .in2(_gnd_net_),
            .in3(N__1544),
            .lcout(\Debounce_Sw1.r_CountZ0Z_2 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_1 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_2 ),
            .clk(N__3081),
            .ce(),
            .sr(N__1802));
    defparam \Debounce_Sw1.r_Count_3_LC_5_5_2 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_3_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_3_LC_5_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_3_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(N__1540),
            .in2(_gnd_net_),
            .in3(N__1526),
            .lcout(\Debounce_Sw1.r_CountZ0Z_3 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_2 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_3 ),
            .clk(N__3081),
            .ce(),
            .sr(N__1802));
    defparam \Debounce_Sw1.r_Count_4_LC_5_5_3 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_4_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_4_LC_5_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_4_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(N__1523),
            .in2(_gnd_net_),
            .in3(N__1511),
            .lcout(\Debounce_Sw1.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_3 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_4 ),
            .clk(N__3081),
            .ce(),
            .sr(N__1802));
    defparam \Debounce_Sw1.r_Count_5_LC_5_5_4 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_5_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_5_LC_5_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_5_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(N__1685),
            .in2(_gnd_net_),
            .in3(N__1673),
            .lcout(\Debounce_Sw1.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_4 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_5 ),
            .clk(N__3081),
            .ce(),
            .sr(N__1802));
    defparam \Debounce_Sw1.r_Count_6_LC_5_5_5 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_6_LC_5_5_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_6_LC_5_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_6_LC_5_5_5  (
            .in0(_gnd_net_),
            .in1(N__2422),
            .in2(_gnd_net_),
            .in3(N__1670),
            .lcout(\Debounce_Sw1.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_5 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_6 ),
            .clk(N__3081),
            .ce(),
            .sr(N__1802));
    defparam \Debounce_Sw1.r_Count_7_LC_5_5_6 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_7_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_7_LC_5_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_7_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(N__2333),
            .in2(_gnd_net_),
            .in3(N__1667),
            .lcout(\Debounce_Sw1.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_6 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_7 ),
            .clk(N__3081),
            .ce(),
            .sr(N__1802));
    defparam \Debounce_Sw1.r_Count_8_LC_5_5_7 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_8_LC_5_5_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_8_LC_5_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_8_LC_5_5_7  (
            .in0(_gnd_net_),
            .in1(N__2443),
            .in2(_gnd_net_),
            .in3(N__1664),
            .lcout(\Debounce_Sw1.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_7 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_8 ),
            .clk(N__3081),
            .ce(),
            .sr(N__1802));
    defparam \Debounce_Sw1.r_Count_9_LC_5_6_0 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_9_LC_5_6_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_9_LC_5_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_9_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(N__2305),
            .in2(_gnd_net_),
            .in3(N__1661),
            .lcout(\Debounce_Sw1.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_5_6_0_),
            .carryout(\Debounce_Sw1.un2_r_count_cry_9 ),
            .clk(N__3079),
            .ce(),
            .sr(N__1801));
    defparam \Debounce_Sw1.r_Count_10_LC_5_6_1 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_10_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_10_LC_5_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_10_LC_5_6_1  (
            .in0(_gnd_net_),
            .in1(N__2284),
            .in2(_gnd_net_),
            .in3(N__1658),
            .lcout(\Debounce_Sw1.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_9 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_10 ),
            .clk(N__3079),
            .ce(),
            .sr(N__1801));
    defparam \Debounce_Sw1.r_Count_11_LC_5_6_2 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_11_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_11_LC_5_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_11_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__2167),
            .in2(_gnd_net_),
            .in3(N__1655),
            .lcout(\Debounce_Sw1.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_10 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_11 ),
            .clk(N__3079),
            .ce(),
            .sr(N__1801));
    defparam \Debounce_Sw1.r_Count_12_LC_5_6_3 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_12_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_12_LC_5_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_12_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(N__2390),
            .in2(_gnd_net_),
            .in3(N__1652),
            .lcout(\Debounce_Sw1.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_11 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_12 ),
            .clk(N__3079),
            .ce(),
            .sr(N__1801));
    defparam \Debounce_Sw1.r_Count_13_LC_5_6_4 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_13_LC_5_6_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_13_LC_5_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_13_LC_5_6_4  (
            .in0(_gnd_net_),
            .in1(N__2213),
            .in2(_gnd_net_),
            .in3(N__1649),
            .lcout(\Debounce_Sw1.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_12 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_13 ),
            .clk(N__3079),
            .ce(),
            .sr(N__1801));
    defparam \Debounce_Sw1.r_Count_14_LC_5_6_5 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_14_LC_5_6_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_14_LC_5_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_14_LC_5_6_5  (
            .in0(_gnd_net_),
            .in1(N__2372),
            .in2(_gnd_net_),
            .in3(N__1814),
            .lcout(\Debounce_Sw1.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_13 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_14 ),
            .clk(N__3079),
            .ce(),
            .sr(N__1801));
    defparam \Debounce_Sw1.r_Count_15_LC_5_6_6 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_15_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_15_LC_5_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_15_LC_5_6_6  (
            .in0(_gnd_net_),
            .in1(N__2353),
            .in2(_gnd_net_),
            .in3(N__1811),
            .lcout(\Debounce_Sw1.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_14 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_15 ),
            .clk(N__3079),
            .ce(),
            .sr(N__1801));
    defparam \Debounce_Sw1.r_Count_16_LC_5_6_7 .C_ON=1'b1;
    defparam \Debounce_Sw1.r_Count_16_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_16_LC_5_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw1.r_Count_16_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(N__2233),
            .in2(_gnd_net_),
            .in3(N__1808),
            .lcout(\Debounce_Sw1.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Debounce_Sw1.un2_r_count_cry_15 ),
            .carryout(\Debounce_Sw1.un2_r_count_cry_16 ),
            .clk(N__3079),
            .ce(),
            .sr(N__1801));
    defparam \Debounce_Sw1.r_Count_17_LC_5_7_0 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_Count_17_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_Count_17_LC_5_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Debounce_Sw1.r_Count_17_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(N__2190),
            .in2(_gnd_net_),
            .in3(N__1805),
            .lcout(\Debounce_Sw1.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3076),
            .ce(),
            .sr(N__1800));
    defparam \Count_And_Toggle.r_Counter_RNIBHPL1_10_LC_5_8_0 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_RNIBHPL1_10_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNIBHPL1_10_LC_5_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Count_And_Toggle.r_Counter_RNIBHPL1_10_LC_5_8_0  (
            .in0(N__1784),
            .in1(N__1769),
            .in2(N__1757),
            .in3(N__1742),
            .lcout(\Count_And_Toggle.un4_i_enable_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_8_LC_5_8_1 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_8_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_8_LC_5_8_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \Count_And_Toggle.r_Counter_8_LC_5_8_1  (
            .in0(N__2048),
            .in1(N__2571),
            .in2(N__2110),
            .in3(N__1730),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3071),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_1_LC_5_8_2 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_1_LC_5_8_2 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_1_LC_5_8_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Count_And_Toggle.r_Counter_1_LC_5_8_2  (
            .in0(N__1858),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1979),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3071),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_0_LC_5_8_3 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_0_LC_5_8_3 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_0_LC_5_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Count_And_Toggle.r_Counter_0_LC_5_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1857),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3071),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNI6J0M1_4_LC_5_8_4 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_RNI6J0M1_4_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNI6J0M1_4_LC_5_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Count_And_Toggle.r_Counter_RNI6J0M1_4_LC_5_8_4  (
            .in0(N__1723),
            .in1(N__1709),
            .in2(N__2132),
            .in3(N__1697),
            .lcout(\Count_And_Toggle.un4_i_enable_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_11_LC_5_8_5 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_11_LC_5_8_5 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_11_LC_5_8_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \Count_And_Toggle.r_Counter_11_LC_5_8_5  (
            .in0(N__2044),
            .in1(N__2569),
            .in2(N__2109),
            .in3(N__2009),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3071),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNIO40M1_1_LC_5_8_6 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_RNIO40M1_1_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNIO40M1_1_LC_5_8_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Count_And_Toggle.r_Counter_RNIO40M1_1_LC_5_8_6  (
            .in0(N__2003),
            .in1(N__1991),
            .in2(N__1955),
            .in3(N__1978),
            .lcout(\Count_And_Toggle.un4_i_enable_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_6_LC_5_8_7 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_6_LC_5_8_7 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_6_LC_5_8_7 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \Count_And_Toggle.r_Counter_6_LC_5_8_7  (
            .in0(N__2100),
            .in1(N__1964),
            .in2(N__2051),
            .in3(N__2570),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3071),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_19_LC_5_9_0 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_19_LC_5_9_0 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_19_LC_5_9_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \Count_And_Toggle.r_Counter_19_LC_5_9_0  (
            .in0(N__2567),
            .in1(N__2042),
            .in2(N__2104),
            .in3(N__1940),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3077),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNI6LNL1_11_LC_5_9_2 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_RNI6LNL1_11_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNI6LNL1_11_LC_5_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Count_And_Toggle.r_Counter_RNI6LNL1_11_LC_5_9_2  (
            .in0(N__1895),
            .in1(N__2456),
            .in2(N__1934),
            .in3(N__1916),
            .lcout(\Count_And_Toggle.un4_i_enable_15 ),
            .ltout(\Count_And_Toggle.un4_i_enable_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_18_LC_5_9_3 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_18_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_18_LC_5_9_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \Count_And_Toggle.r_Counter_18_LC_5_9_3  (
            .in0(N__2090),
            .in1(N__2566),
            .in2(N__1904),
            .in3(N__1901),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3077),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNIMOB81_15_LC_5_9_4 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_RNIMOB81_15_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNIMOB81_15_LC_5_9_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Count_And_Toggle.r_Counter_RNIMOB81_15_LC_5_9_4  (
            .in0(N__1883),
            .in1(N__1871),
            .in2(_gnd_net_),
            .in3(N__1856),
            .lcout(),
            .ltout(\Count_And_Toggle.un4_i_enable_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_RNIV16A6_10_LC_5_9_5 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_RNIV16A6_10_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \Count_And_Toggle.r_Counter_RNIV16A6_10_LC_5_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Count_And_Toggle.r_Counter_RNIV16A6_10_LC_5_9_5  (
            .in0(N__1835),
            .in1(N__1829),
            .in2(N__1823),
            .in3(N__1820),
            .lcout(\Count_And_Toggle.un4_i_enable_20 ),
            .ltout(\Count_And_Toggle.un4_i_enable_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_14_LC_5_9_6 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_14_LC_5_9_6 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_14_LC_5_9_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \Count_And_Toggle.r_Counter_14_LC_5_9_6  (
            .in0(N__2086),
            .in1(N__2041),
            .in2(N__2465),
            .in3(N__2462),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3077),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.r_State_RNO_0_LC_6_5_5 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_State_RNO_0_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw1.r_State_RNO_0_LC_6_5_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Debounce_Sw1.r_State_RNO_0_LC_6_5_5  (
            .in0(N__2444),
            .in1(N__2147),
            .in2(N__2426),
            .in3(N__2405),
            .lcout(\Debounce_Sw1.un9_r_count_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.r_State_RNO_3_LC_6_6_4 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_State_RNO_3_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw1.r_State_RNO_3_LC_6_6_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_Sw1.r_State_RNO_3_LC_6_6_4  (
            .in0(N__2389),
            .in1(N__2371),
            .in2(N__2354),
            .in3(N__2332),
            .lcout(),
            .ltout(\Debounce_Sw1.un9_r_count_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.r_State_RNO_1_LC_6_6_5 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_State_RNO_1_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw1.r_State_RNO_1_LC_6_6_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Debounce_Sw1.r_State_RNO_1_LC_6_6_5  (
            .in0(N__2315),
            .in1(N__2306),
            .in2(N__2288),
            .in3(N__2285),
            .lcout(),
            .ltout(\Debounce_Sw1.un9_r_count_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.r_State_LC_6_6_6 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_State_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw1.r_State_LC_6_6_6 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Debounce_Sw1.r_State_LC_6_6_6  (
            .in0(N__2267),
            .in1(N__2254),
            .in2(N__2237),
            .in3(N__2973),
            .lcout(w_Switch_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3083),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw1.r_State_RNO_2_LC_6_6_7 .C_ON=1'b0;
    defparam \Debounce_Sw1.r_State_RNO_2_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw1.r_State_RNO_2_LC_6_6_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Debounce_Sw1.r_State_RNO_2_LC_6_6_7  (
            .in0(N__2232),
            .in1(N__2212),
            .in2(N__2194),
            .in3(N__2166),
            .lcout(\Debounce_Sw1.un9_r_count_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.r_Counter_9_LC_6_8_5 .C_ON=1'b0;
    defparam \Count_And_Toggle.r_Counter_9_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.r_Counter_9_LC_6_8_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \Count_And_Toggle.r_Counter_9_LC_6_8_5  (
            .in0(N__2050),
            .in1(N__2573),
            .in2(N__2114),
            .in3(N__2141),
            .lcout(\Count_And_Toggle.r_CounterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3074),
            .ce(),
            .sr(_gnd_net_));
    defparam \Count_And_Toggle.o_Toggle_LC_6_9_0 .C_ON=1'b0;
    defparam \Count_And_Toggle.o_Toggle_LC_6_9_0 .SEQ_MODE=4'b1000;
    defparam \Count_And_Toggle.o_Toggle_LC_6_9_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \Count_And_Toggle.o_Toggle_LC_6_9_0  (
            .in0(N__2105),
            .in1(N__2043),
            .in2(N__2935),
            .in3(N__2568),
            .lcout(w_Toggle),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3080),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw2.r_State_e_0_LC_6_10_1 .C_ON=1'b0;
    defparam \Debounce_Sw2.r_State_e_0_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_State_e_0_LC_6_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Debounce_Sw2.r_State_e_0_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2524),
            .lcout(w_Switch_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3082),
            .ce(N__2474),
            .sr(_gnd_net_));
    defparam \Debounce_Sw2.r_Count_1_LC_7_8_0 .C_ON=1'b0;
    defparam \Debounce_Sw2.r_Count_1_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_1_LC_7_8_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Debounce_Sw2.r_Count_1_LC_7_8_0  (
            .in0(N__2684),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2662),
            .lcout(\Debounce_Sw2.r_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3078),
            .ce(),
            .sr(N__3028));
    defparam \Debounce_Sw2.r_Count_0_LC_7_8_7 .C_ON=1'b0;
    defparam \Debounce_Sw2.r_Count_0_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_0_LC_7_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Debounce_Sw2.r_Count_0_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2683),
            .lcout(\Debounce_Sw2.r_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3078),
            .ce(),
            .sr(N__3028));
    defparam \Debounce_Sw2.r_Count_RNIV5631_4_LC_7_9_0 .C_ON=1'b0;
    defparam \Debounce_Sw2.r_Count_RNIV5631_4_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw2.r_Count_RNIV5631_4_LC_7_9_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Debounce_Sw2.r_Count_RNIV5631_4_LC_7_9_0  (
            .in0(N__2591),
            .in1(N__2605),
            .in2(_gnd_net_),
            .in3(N__2875),
            .lcout(\Debounce_Sw2.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw2.r_Count_RNI64TE1_1_LC_7_9_2 .C_ON=1'b0;
    defparam \Debounce_Sw2.r_Count_RNI64TE1_1_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw2.r_Count_RNI64TE1_1_LC_7_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_Sw2.r_Count_RNI64TE1_1_LC_7_9_2  (
            .in0(N__2620),
            .in1(N__2658),
            .in2(N__2642),
            .in3(N__2681),
            .lcout(\Debounce_Sw2.un9_r_count_10 ),
            .ltout(\Debounce_Sw2.un9_r_count_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw2.r_Count_RNISOQT2_7_LC_7_9_3 .C_ON=1'b0;
    defparam \Debounce_Sw2.r_Count_RNISOQT2_7_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw2.r_Count_RNISOQT2_7_LC_7_9_3 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \Debounce_Sw2.r_Count_RNISOQT2_7_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(N__2856),
            .in2(N__2534),
            .in3(N__2719),
            .lcout(),
            .ltout(\Debounce_Sw2.N_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw2.r_Count_RNINN314_12_LC_7_9_4 .C_ON=1'b0;
    defparam \Debounce_Sw2.r_Count_RNINN314_12_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw2.r_Count_RNINN314_12_LC_7_9_4 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \Debounce_Sw2.r_Count_RNINN314_12_LC_7_9_4  (
            .in0(N__2772),
            .in1(N__2754),
            .in2(N__2531),
            .in3(N__2692),
            .lcout(),
            .ltout(\Debounce_Sw2.N_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw2.r_State_e_0_RNIK82U4_LC_7_9_5 .C_ON=1'b0;
    defparam \Debounce_Sw2.r_State_e_0_RNIK82U4_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw2.r_State_e_0_RNIK82U4_LC_7_9_5 .LUT_INIT=16'b1110101011010101;
    LogicCell40 \Debounce_Sw2.r_State_e_0_RNIK82U4_LC_7_9_5  (
            .in0(N__2528),
            .in1(N__2701),
            .in2(N__2498),
            .in3(N__2893),
            .lcout(\Debounce_Sw2.N_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw2.r_State_e_0_RNO_LC_7_9_6 .C_ON=1'b0;
    defparam \Debounce_Sw2.r_State_e_0_RNO_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw2.r_State_e_0_RNO_LC_7_9_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Debounce_Sw2.r_State_e_0_RNO_LC_7_9_6  (
            .in0(N__2702),
            .in1(N__2708),
            .in2(N__2483),
            .in3(N__2693),
            .lcout(\Debounce_Sw2.r_State_e_0_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw2.r_State_e_0_RNO_0_LC_7_9_7 .C_ON=1'b0;
    defparam \Debounce_Sw2.r_State_e_0_RNO_0_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw2.r_State_e_0_RNO_0_LC_7_9_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Debounce_Sw2.r_State_e_0_RNO_0_LC_7_9_7  (
            .in0(N__2720),
            .in1(N__2773),
            .in2(N__2861),
            .in3(N__2755),
            .lcout(\Debounce_Sw2.un9_r_count_0_a3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw2.r_Count_RNIQEQB_17_LC_7_10_0 .C_ON=1'b0;
    defparam \Debounce_Sw2.r_Count_RNIQEQB_17_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw2.r_Count_RNIQEQB_17_LC_7_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_Sw2.r_Count_RNIQEQB_17_LC_7_10_0  (
            .in0(N__3121),
            .in1(N__3136),
            .in2(N__3104),
            .in3(N__2734),
            .lcout(\Debounce_Sw2.N_22_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw2.r_Count_RNIKTBT_10_LC_7_10_5 .C_ON=1'b0;
    defparam \Debounce_Sw2.r_Count_RNIKTBT_10_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw2.r_Count_RNIKTBT_10_LC_7_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Debounce_Sw2.r_Count_RNIKTBT_10_LC_7_10_5  (
            .in0(N__2806),
            .in1(N__2821),
            .in2(N__2792),
            .in3(N__2836),
            .lcout(\Debounce_Sw2.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw2.un2_r_count_cry_1_c_LC_8_9_0 .C_ON=1'b1;
    defparam \Debounce_Sw2.un2_r_count_cry_1_c_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_Sw2.un2_r_count_cry_1_c_LC_8_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Debounce_Sw2.un2_r_count_cry_1_c_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__2682),
            .in2(N__2663),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\Debounce_Sw2.un2_r_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_Sw2.r_Count_2_LC_8_9_1 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_2_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_2_LC_8_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_2_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__2638),
            .in2(_gnd_net_),
            .in3(N__2624),
            .lcout(\Debounce_Sw2.r_CountZ0Z_2 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_1 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_2 ),
            .clk(N__3084),
            .ce(),
            .sr(N__3029));
    defparam \Debounce_Sw2.r_Count_3_LC_8_9_2 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_3_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_3_LC_8_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_3_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__2621),
            .in2(_gnd_net_),
            .in3(N__2609),
            .lcout(\Debounce_Sw2.r_CountZ0Z_3 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_2 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_3 ),
            .clk(N__3084),
            .ce(),
            .sr(N__3029));
    defparam \Debounce_Sw2.r_Count_4_LC_8_9_3 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_4_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_4_LC_8_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_4_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__2606),
            .in2(_gnd_net_),
            .in3(N__2594),
            .lcout(\Debounce_Sw2.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_3 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_4 ),
            .clk(N__3084),
            .ce(),
            .sr(N__3029));
    defparam \Debounce_Sw2.r_Count_5_LC_8_9_4 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_5_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_5_LC_8_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_5_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__2590),
            .in2(_gnd_net_),
            .in3(N__2576),
            .lcout(\Debounce_Sw2.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_4 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_5 ),
            .clk(N__3084),
            .ce(),
            .sr(N__3029));
    defparam \Debounce_Sw2.r_Count_6_LC_8_9_5 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_6_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_6_LC_8_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_6_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__2876),
            .in2(_gnd_net_),
            .in3(N__2864),
            .lcout(\Debounce_Sw2.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_5 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_6 ),
            .clk(N__3084),
            .ce(),
            .sr(N__3029));
    defparam \Debounce_Sw2.r_Count_7_LC_8_9_6 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_7_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_7_LC_8_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_7_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__2860),
            .in2(_gnd_net_),
            .in3(N__2840),
            .lcout(\Debounce_Sw2.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_6 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_7 ),
            .clk(N__3084),
            .ce(),
            .sr(N__3029));
    defparam \Debounce_Sw2.r_Count_8_LC_8_9_7 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_8_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_8_LC_8_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_8_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__2837),
            .in2(_gnd_net_),
            .in3(N__2825),
            .lcout(\Debounce_Sw2.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_7 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_8 ),
            .clk(N__3084),
            .ce(),
            .sr(N__3029));
    defparam \Debounce_Sw2.r_Count_9_LC_8_10_0 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_9_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_9_LC_8_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_9_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__2822),
            .in2(_gnd_net_),
            .in3(N__2810),
            .lcout(\Debounce_Sw2.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\Debounce_Sw2.un2_r_count_cry_9 ),
            .clk(N__3085),
            .ce(),
            .sr(N__3027));
    defparam \Debounce_Sw2.r_Count_10_LC_8_10_1 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_10_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_10_LC_8_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_10_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__2807),
            .in2(_gnd_net_),
            .in3(N__2795),
            .lcout(\Debounce_Sw2.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_9 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_10 ),
            .clk(N__3085),
            .ce(),
            .sr(N__3027));
    defparam \Debounce_Sw2.r_Count_11_LC_8_10_2 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_11_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_11_LC_8_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_11_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__2791),
            .in2(_gnd_net_),
            .in3(N__2777),
            .lcout(\Debounce_Sw2.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_10 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_11 ),
            .clk(N__3085),
            .ce(),
            .sr(N__3027));
    defparam \Debounce_Sw2.r_Count_12_LC_8_10_3 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_12_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_12_LC_8_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_12_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__2774),
            .in2(_gnd_net_),
            .in3(N__2759),
            .lcout(\Debounce_Sw2.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_11 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_12 ),
            .clk(N__3085),
            .ce(),
            .sr(N__3027));
    defparam \Debounce_Sw2.r_Count_13_LC_8_10_4 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_13_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_13_LC_8_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_13_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__2756),
            .in2(_gnd_net_),
            .in3(N__2738),
            .lcout(\Debounce_Sw2.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_12 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_13 ),
            .clk(N__3085),
            .ce(),
            .sr(N__3027));
    defparam \Debounce_Sw2.r_Count_14_LC_8_10_5 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_14_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_14_LC_8_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_14_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__2735),
            .in2(_gnd_net_),
            .in3(N__2723),
            .lcout(\Debounce_Sw2.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_13 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_14 ),
            .clk(N__3085),
            .ce(),
            .sr(N__3027));
    defparam \Debounce_Sw2.r_Count_15_LC_8_10_6 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_15_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_15_LC_8_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_15_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__3137),
            .in2(_gnd_net_),
            .in3(N__3125),
            .lcout(\Debounce_Sw2.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_14 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_15 ),
            .clk(N__3085),
            .ce(),
            .sr(N__3027));
    defparam \Debounce_Sw2.r_Count_16_LC_8_10_7 .C_ON=1'b1;
    defparam \Debounce_Sw2.r_Count_16_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_16_LC_8_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_Sw2.r_Count_16_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(N__3122),
            .in2(_gnd_net_),
            .in3(N__3110),
            .lcout(\Debounce_Sw2.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Debounce_Sw2.un2_r_count_cry_15 ),
            .carryout(\Debounce_Sw2.un2_r_count_cry_16 ),
            .clk(N__3085),
            .ce(),
            .sr(N__3027));
    defparam \Debounce_Sw2.r_Count_17_LC_8_11_0 .C_ON=1'b0;
    defparam \Debounce_Sw2.r_Count_17_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_Sw2.r_Count_17_LC_8_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Debounce_Sw2.r_Count_17_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__3100),
            .in2(_gnd_net_),
            .in3(N__3107),
            .lcout(\Debounce_Sw2.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3086),
            .ce(),
            .sr(N__3026));
    defparam \Demux.o_Data2_0_a3_LC_12_7_0 .C_ON=1'b0;
    defparam \Demux.o_Data2_0_a3_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \Demux.o_Data2_0_a3_LC_12_7_0 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \Demux.o_Data2_0_a3_LC_12_7_0  (
            .in0(N__2953),
            .in1(_gnd_net_),
            .in2(N__2918),
            .in3(N__2991),
            .lcout(o_LED_2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Demux.o_Data3_0_a3_LC_12_7_1 .C_ON=1'b0;
    defparam \Demux.o_Data3_0_a3_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \Demux.o_Data3_0_a3_LC_12_7_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Demux.o_Data3_0_a3_LC_12_7_1  (
            .in0(N__2992),
            .in1(N__2954),
            .in2(_gnd_net_),
            .in3(N__2917),
            .lcout(o_LED_3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Demux.o_Data1_0_a3_LC_12_7_7 .C_ON=1'b0;
    defparam \Demux.o_Data1_0_a3_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \Demux.o_Data1_0_a3_LC_12_7_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \Demux.o_Data1_0_a3_LC_12_7_7  (
            .in0(N__2990),
            .in1(N__2952),
            .in2(_gnd_net_),
            .in3(N__2913),
            .lcout(o_LED_1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Demux.o_Data4_0_a3_LC_12_8_1 .C_ON=1'b0;
    defparam \Demux.o_Data4_0_a3_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \Demux.o_Data4_0_a3_LC_12_8_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Demux.o_Data4_0_a3_LC_12_8_1  (
            .in0(N__2993),
            .in1(N__2951),
            .in2(_gnd_net_),
            .in3(N__2912),
            .lcout(o_LED_4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // Demux_Toggle_TOP
